module rom_data (
    input wire [15:0] addr,
    output reg [2:0] data
);

    reg [2:0] rom_memory [0:52799];  // 240 * 220 = 52800

    initial begin
        rom_memory[0] = 3'b110;
        rom_memory[1] = 3'b110;
        rom_memory[2] = 3'b110;
        rom_memory[3] = 3'b110;
        rom_memory[4] = 3'b110;
        rom_memory[5] = 3'b110;
        rom_memory[6] = 3'b110;
        rom_memory[7] = 3'b110;
        rom_memory[8] = 3'b110;
        rom_memory[9] = 3'b110;
        rom_memory[10] = 3'b110;
        rom_memory[11] = 3'b110;
        rom_memory[12] = 3'b110;
        rom_memory[13] = 3'b110;
        rom_memory[14] = 3'b110;
        rom_memory[15] = 3'b110;
        rom_memory[16] = 3'b110;
        rom_memory[17] = 3'b110;
        rom_memory[18] = 3'b110;
        rom_memory[19] = 3'b110;
        rom_memory[20] = 3'b110;
        rom_memory[21] = 3'b110;
        rom_memory[22] = 3'b110;
        rom_memory[23] = 3'b110;
        rom_memory[24] = 3'b110;
        rom_memory[25] = 3'b110;
        rom_memory[26] = 3'b110;
        rom_memory[27] = 3'b110;
        rom_memory[28] = 3'b110;
        rom_memory[29] = 3'b110;
        rom_memory[30] = 3'b110;
        rom_memory[31] = 3'b110;
        rom_memory[32] = 3'b110;
        rom_memory[33] = 3'b110;
        rom_memory[34] = 3'b110;
        rom_memory[35] = 3'b110;
        rom_memory[36] = 3'b110;
        rom_memory[37] = 3'b110;
        rom_memory[38] = 3'b110;
        rom_memory[39] = 3'b110;
        rom_memory[40] = 3'b110;
        rom_memory[41] = 3'b110;
        rom_memory[42] = 3'b110;
        rom_memory[43] = 3'b110;
        rom_memory[44] = 3'b110;
        rom_memory[45] = 3'b110;
        rom_memory[46] = 3'b110;
        rom_memory[47] = 3'b110;
        rom_memory[48] = 3'b110;
        rom_memory[49] = 3'b110;
        rom_memory[50] = 3'b110;
        rom_memory[51] = 3'b110;
        rom_memory[52] = 3'b110;
        rom_memory[53] = 3'b110;
        rom_memory[54] = 3'b110;
        rom_memory[55] = 3'b110;
        rom_memory[56] = 3'b110;
        rom_memory[57] = 3'b110;
        rom_memory[58] = 3'b110;
        rom_memory[59] = 3'b110;
        rom_memory[60] = 3'b110;
        rom_memory[61] = 3'b110;
        rom_memory[62] = 3'b110;
        rom_memory[63] = 3'b110;
        rom_memory[64] = 3'b110;
        rom_memory[65] = 3'b110;
        rom_memory[66] = 3'b110;
        rom_memory[67] = 3'b110;
        rom_memory[68] = 3'b110;
        rom_memory[69] = 3'b110;
        rom_memory[70] = 3'b110;
        rom_memory[71] = 3'b110;
        rom_memory[72] = 3'b110;
        rom_memory[73] = 3'b110;
        rom_memory[74] = 3'b110;
        rom_memory[75] = 3'b110;
        rom_memory[76] = 3'b110;
        rom_memory[77] = 3'b110;
        rom_memory[78] = 3'b110;
        rom_memory[79] = 3'b110;
        rom_memory[80] = 3'b110;
        rom_memory[81] = 3'b110;
        rom_memory[82] = 3'b110;
        rom_memory[83] = 3'b110;
        rom_memory[84] = 3'b110;
        rom_memory[85] = 3'b110;
        rom_memory[86] = 3'b110;
        rom_memory[87] = 3'b110;
        rom_memory[88] = 3'b110;
        rom_memory[89] = 3'b110;
        rom_memory[90] = 3'b110;
        rom_memory[91] = 3'b110;
        rom_memory[92] = 3'b110;
        rom_memory[93] = 3'b110;
        rom_memory[94] = 3'b110;
        rom_memory[95] = 3'b110;
        rom_memory[96] = 3'b110;
        rom_memory[97] = 3'b110;
        rom_memory[98] = 3'b110;
        rom_memory[99] = 3'b110;
        rom_memory[100] = 3'b110;
        rom_memory[101] = 3'b110;
        rom_memory[102] = 3'b110;
        rom_memory[103] = 3'b110;
        rom_memory[104] = 3'b110;
        rom_memory[105] = 3'b110;
        rom_memory[106] = 3'b110;
        rom_memory[107] = 3'b110;
        rom_memory[108] = 3'b110;
        rom_memory[109] = 3'b110;
        rom_memory[110] = 3'b110;
        rom_memory[111] = 3'b110;
        rom_memory[112] = 3'b110;
        rom_memory[113] = 3'b110;
        rom_memory[114] = 3'b110;
        rom_memory[115] = 3'b110;
        rom_memory[116] = 3'b110;
        rom_memory[117] = 3'b110;
        rom_memory[118] = 3'b110;
        rom_memory[119] = 3'b110;
        rom_memory[120] = 3'b110;
        rom_memory[121] = 3'b110;
        rom_memory[122] = 3'b110;
        rom_memory[123] = 3'b110;
        rom_memory[124] = 3'b110;
        rom_memory[125] = 3'b110;
        rom_memory[126] = 3'b110;
        rom_memory[127] = 3'b110;
        rom_memory[128] = 3'b110;
        rom_memory[129] = 3'b110;
        rom_memory[130] = 3'b110;
        rom_memory[131] = 3'b110;
        rom_memory[132] = 3'b110;
        rom_memory[133] = 3'b110;
        rom_memory[134] = 3'b110;
        rom_memory[135] = 3'b110;
        rom_memory[136] = 3'b110;
        rom_memory[137] = 3'b110;
        rom_memory[138] = 3'b110;
        rom_memory[139] = 3'b110;
        rom_memory[140] = 3'b110;
        rom_memory[141] = 3'b110;
        rom_memory[142] = 3'b110;
        rom_memory[143] = 3'b110;
        rom_memory[144] = 3'b110;
        rom_memory[145] = 3'b110;
        rom_memory[146] = 3'b110;
        rom_memory[147] = 3'b110;
        rom_memory[148] = 3'b110;
        rom_memory[149] = 3'b110;
        rom_memory[150] = 3'b110;
        rom_memory[151] = 3'b110;
        rom_memory[152] = 3'b110;
        rom_memory[153] = 3'b110;
        rom_memory[154] = 3'b110;
        rom_memory[155] = 3'b110;
        rom_memory[156] = 3'b110;
        rom_memory[157] = 3'b110;
        rom_memory[158] = 3'b110;
        rom_memory[159] = 3'b100;
        rom_memory[160] = 3'b100;
        rom_memory[161] = 3'b100;
        rom_memory[162] = 3'b100;
        rom_memory[163] = 3'b100;
        rom_memory[164] = 3'b100;
        rom_memory[165] = 3'b100;
        rom_memory[166] = 3'b100;
        rom_memory[167] = 3'b100;
        rom_memory[168] = 3'b100;
        rom_memory[169] = 3'b100;
        rom_memory[170] = 3'b100;
        rom_memory[171] = 3'b100;
        rom_memory[172] = 3'b100;
        rom_memory[173] = 3'b100;
        rom_memory[174] = 3'b100;
        rom_memory[175] = 3'b100;
        rom_memory[176] = 3'b100;
        rom_memory[177] = 3'b100;
        rom_memory[178] = 3'b100;
        rom_memory[179] = 3'b100;
        rom_memory[180] = 3'b100;
        rom_memory[181] = 3'b100;
        rom_memory[182] = 3'b100;
        rom_memory[183] = 3'b100;
        rom_memory[184] = 3'b100;
        rom_memory[185] = 3'b100;
        rom_memory[186] = 3'b100;
        rom_memory[187] = 3'b100;
        rom_memory[188] = 3'b100;
        rom_memory[189] = 3'b100;
        rom_memory[190] = 3'b100;
        rom_memory[191] = 3'b100;
        rom_memory[192] = 3'b100;
        rom_memory[193] = 3'b100;
        rom_memory[194] = 3'b100;
        rom_memory[195] = 3'b100;
        rom_memory[196] = 3'b100;
        rom_memory[197] = 3'b100;
        rom_memory[198] = 3'b100;
        rom_memory[199] = 3'b100;
        rom_memory[200] = 3'b100;
        rom_memory[201] = 3'b100;
        rom_memory[202] = 3'b100;
        rom_memory[203] = 3'b100;
        rom_memory[204] = 3'b100;
        rom_memory[205] = 3'b100;
        rom_memory[206] = 3'b100;
        rom_memory[207] = 3'b100;
        rom_memory[208] = 3'b100;
        rom_memory[209] = 3'b100;
        rom_memory[210] = 3'b100;
        rom_memory[211] = 3'b100;
        rom_memory[212] = 3'b100;
        rom_memory[213] = 3'b100;
        rom_memory[214] = 3'b100;
        rom_memory[215] = 3'b100;
        rom_memory[216] = 3'b100;
        rom_memory[217] = 3'b100;
        rom_memory[218] = 3'b100;
        rom_memory[219] = 3'b100;
        rom_memory[220] = 3'b100;
        rom_memory[221] = 3'b100;
        rom_memory[222] = 3'b100;
        rom_memory[223] = 3'b100;
        rom_memory[224] = 3'b100;
        rom_memory[225] = 3'b100;
        rom_memory[226] = 3'b100;
        rom_memory[227] = 3'b100;
        rom_memory[228] = 3'b100;
        rom_memory[229] = 3'b100;
        rom_memory[230] = 3'b100;
        rom_memory[231] = 3'b100;
        rom_memory[232] = 3'b100;
        rom_memory[233] = 3'b100;
        rom_memory[234] = 3'b100;
        rom_memory[235] = 3'b100;
        rom_memory[236] = 3'b100;
        rom_memory[237] = 3'b100;
        rom_memory[238] = 3'b100;
        rom_memory[239] = 3'b100;
        rom_memory[240] = 3'b110;
        rom_memory[241] = 3'b110;
        rom_memory[242] = 3'b110;
        rom_memory[243] = 3'b110;
        rom_memory[244] = 3'b110;
        rom_memory[245] = 3'b110;
        rom_memory[246] = 3'b110;
        rom_memory[247] = 3'b110;
        rom_memory[248] = 3'b110;
        rom_memory[249] = 3'b110;
        rom_memory[250] = 3'b110;
        rom_memory[251] = 3'b110;
        rom_memory[252] = 3'b110;
        rom_memory[253] = 3'b110;
        rom_memory[254] = 3'b110;
        rom_memory[255] = 3'b110;
        rom_memory[256] = 3'b110;
        rom_memory[257] = 3'b110;
        rom_memory[258] = 3'b110;
        rom_memory[259] = 3'b110;
        rom_memory[260] = 3'b110;
        rom_memory[261] = 3'b110;
        rom_memory[262] = 3'b110;
        rom_memory[263] = 3'b110;
        rom_memory[264] = 3'b110;
        rom_memory[265] = 3'b110;
        rom_memory[266] = 3'b110;
        rom_memory[267] = 3'b110;
        rom_memory[268] = 3'b110;
        rom_memory[269] = 3'b110;
        rom_memory[270] = 3'b110;
        rom_memory[271] = 3'b110;
        rom_memory[272] = 3'b110;
        rom_memory[273] = 3'b110;
        rom_memory[274] = 3'b110;
        rom_memory[275] = 3'b110;
        rom_memory[276] = 3'b110;
        rom_memory[277] = 3'b110;
        rom_memory[278] = 3'b110;
        rom_memory[279] = 3'b110;
        rom_memory[280] = 3'b110;
        rom_memory[281] = 3'b110;
        rom_memory[282] = 3'b110;
        rom_memory[283] = 3'b110;
        rom_memory[284] = 3'b110;
        rom_memory[285] = 3'b110;
        rom_memory[286] = 3'b110;
        rom_memory[287] = 3'b110;
        rom_memory[288] = 3'b110;
        rom_memory[289] = 3'b110;
        rom_memory[290] = 3'b110;
        rom_memory[291] = 3'b110;
        rom_memory[292] = 3'b110;
        rom_memory[293] = 3'b110;
        rom_memory[294] = 3'b110;
        rom_memory[295] = 3'b110;
        rom_memory[296] = 3'b110;
        rom_memory[297] = 3'b110;
        rom_memory[298] = 3'b110;
        rom_memory[299] = 3'b110;
        rom_memory[300] = 3'b110;
        rom_memory[301] = 3'b110;
        rom_memory[302] = 3'b110;
        rom_memory[303] = 3'b110;
        rom_memory[304] = 3'b110;
        rom_memory[305] = 3'b110;
        rom_memory[306] = 3'b110;
        rom_memory[307] = 3'b110;
        rom_memory[308] = 3'b110;
        rom_memory[309] = 3'b110;
        rom_memory[310] = 3'b110;
        rom_memory[311] = 3'b110;
        rom_memory[312] = 3'b110;
        rom_memory[313] = 3'b110;
        rom_memory[314] = 3'b110;
        rom_memory[315] = 3'b110;
        rom_memory[316] = 3'b110;
        rom_memory[317] = 3'b110;
        rom_memory[318] = 3'b110;
        rom_memory[319] = 3'b110;
        rom_memory[320] = 3'b110;
        rom_memory[321] = 3'b110;
        rom_memory[322] = 3'b110;
        rom_memory[323] = 3'b110;
        rom_memory[324] = 3'b110;
        rom_memory[325] = 3'b110;
        rom_memory[326] = 3'b110;
        rom_memory[327] = 3'b110;
        rom_memory[328] = 3'b110;
        rom_memory[329] = 3'b110;
        rom_memory[330] = 3'b110;
        rom_memory[331] = 3'b110;
        rom_memory[332] = 3'b110;
        rom_memory[333] = 3'b110;
        rom_memory[334] = 3'b110;
        rom_memory[335] = 3'b110;
        rom_memory[336] = 3'b110;
        rom_memory[337] = 3'b110;
        rom_memory[338] = 3'b110;
        rom_memory[339] = 3'b110;
        rom_memory[340] = 3'b110;
        rom_memory[341] = 3'b110;
        rom_memory[342] = 3'b110;
        rom_memory[343] = 3'b110;
        rom_memory[344] = 3'b110;
        rom_memory[345] = 3'b110;
        rom_memory[346] = 3'b110;
        rom_memory[347] = 3'b110;
        rom_memory[348] = 3'b110;
        rom_memory[349] = 3'b110;
        rom_memory[350] = 3'b110;
        rom_memory[351] = 3'b110;
        rom_memory[352] = 3'b110;
        rom_memory[353] = 3'b110;
        rom_memory[354] = 3'b110;
        rom_memory[355] = 3'b110;
        rom_memory[356] = 3'b110;
        rom_memory[357] = 3'b110;
        rom_memory[358] = 3'b110;
        rom_memory[359] = 3'b110;
        rom_memory[360] = 3'b110;
        rom_memory[361] = 3'b110;
        rom_memory[362] = 3'b110;
        rom_memory[363] = 3'b110;
        rom_memory[364] = 3'b110;
        rom_memory[365] = 3'b110;
        rom_memory[366] = 3'b110;
        rom_memory[367] = 3'b110;
        rom_memory[368] = 3'b110;
        rom_memory[369] = 3'b110;
        rom_memory[370] = 3'b110;
        rom_memory[371] = 3'b110;
        rom_memory[372] = 3'b110;
        rom_memory[373] = 3'b110;
        rom_memory[374] = 3'b110;
        rom_memory[375] = 3'b110;
        rom_memory[376] = 3'b110;
        rom_memory[377] = 3'b110;
        rom_memory[378] = 3'b110;
        rom_memory[379] = 3'b110;
        rom_memory[380] = 3'b110;
        rom_memory[381] = 3'b110;
        rom_memory[382] = 3'b110;
        rom_memory[383] = 3'b110;
        rom_memory[384] = 3'b110;
        rom_memory[385] = 3'b110;
        rom_memory[386] = 3'b110;
        rom_memory[387] = 3'b110;
        rom_memory[388] = 3'b110;
        rom_memory[389] = 3'b110;
        rom_memory[390] = 3'b110;
        rom_memory[391] = 3'b110;
        rom_memory[392] = 3'b110;
        rom_memory[393] = 3'b110;
        rom_memory[394] = 3'b110;
        rom_memory[395] = 3'b110;
        rom_memory[396] = 3'b110;
        rom_memory[397] = 3'b110;
        rom_memory[398] = 3'b110;
        rom_memory[399] = 3'b100;
        rom_memory[400] = 3'b100;
        rom_memory[401] = 3'b100;
        rom_memory[402] = 3'b100;
        rom_memory[403] = 3'b100;
        rom_memory[404] = 3'b100;
        rom_memory[405] = 3'b100;
        rom_memory[406] = 3'b100;
        rom_memory[407] = 3'b100;
        rom_memory[408] = 3'b100;
        rom_memory[409] = 3'b100;
        rom_memory[410] = 3'b100;
        rom_memory[411] = 3'b100;
        rom_memory[412] = 3'b100;
        rom_memory[413] = 3'b100;
        rom_memory[414] = 3'b100;
        rom_memory[415] = 3'b100;
        rom_memory[416] = 3'b100;
        rom_memory[417] = 3'b100;
        rom_memory[418] = 3'b100;
        rom_memory[419] = 3'b100;
        rom_memory[420] = 3'b100;
        rom_memory[421] = 3'b100;
        rom_memory[422] = 3'b100;
        rom_memory[423] = 3'b100;
        rom_memory[424] = 3'b100;
        rom_memory[425] = 3'b100;
        rom_memory[426] = 3'b100;
        rom_memory[427] = 3'b100;
        rom_memory[428] = 3'b100;
        rom_memory[429] = 3'b100;
        rom_memory[430] = 3'b100;
        rom_memory[431] = 3'b100;
        rom_memory[432] = 3'b100;
        rom_memory[433] = 3'b100;
        rom_memory[434] = 3'b100;
        rom_memory[435] = 3'b100;
        rom_memory[436] = 3'b100;
        rom_memory[437] = 3'b100;
        rom_memory[438] = 3'b100;
        rom_memory[439] = 3'b100;
        rom_memory[440] = 3'b100;
        rom_memory[441] = 3'b100;
        rom_memory[442] = 3'b100;
        rom_memory[443] = 3'b100;
        rom_memory[444] = 3'b100;
        rom_memory[445] = 3'b100;
        rom_memory[446] = 3'b100;
        rom_memory[447] = 3'b100;
        rom_memory[448] = 3'b100;
        rom_memory[449] = 3'b100;
        rom_memory[450] = 3'b100;
        rom_memory[451] = 3'b100;
        rom_memory[452] = 3'b100;
        rom_memory[453] = 3'b100;
        rom_memory[454] = 3'b100;
        rom_memory[455] = 3'b100;
        rom_memory[456] = 3'b100;
        rom_memory[457] = 3'b100;
        rom_memory[458] = 3'b100;
        rom_memory[459] = 3'b100;
        rom_memory[460] = 3'b100;
        rom_memory[461] = 3'b100;
        rom_memory[462] = 3'b100;
        rom_memory[463] = 3'b100;
        rom_memory[464] = 3'b100;
        rom_memory[465] = 3'b100;
        rom_memory[466] = 3'b100;
        rom_memory[467] = 3'b100;
        rom_memory[468] = 3'b100;
        rom_memory[469] = 3'b100;
        rom_memory[470] = 3'b100;
        rom_memory[471] = 3'b100;
        rom_memory[472] = 3'b100;
        rom_memory[473] = 3'b100;
        rom_memory[474] = 3'b100;
        rom_memory[475] = 3'b100;
        rom_memory[476] = 3'b100;
        rom_memory[477] = 3'b100;
        rom_memory[478] = 3'b100;
        rom_memory[479] = 3'b100;
        rom_memory[480] = 3'b110;
        rom_memory[481] = 3'b110;
        rom_memory[482] = 3'b110;
        rom_memory[483] = 3'b110;
        rom_memory[484] = 3'b110;
        rom_memory[485] = 3'b110;
        rom_memory[486] = 3'b110;
        rom_memory[487] = 3'b110;
        rom_memory[488] = 3'b110;
        rom_memory[489] = 3'b110;
        rom_memory[490] = 3'b110;
        rom_memory[491] = 3'b110;
        rom_memory[492] = 3'b110;
        rom_memory[493] = 3'b110;
        rom_memory[494] = 3'b110;
        rom_memory[495] = 3'b110;
        rom_memory[496] = 3'b110;
        rom_memory[497] = 3'b110;
        rom_memory[498] = 3'b110;
        rom_memory[499] = 3'b110;
        rom_memory[500] = 3'b110;
        rom_memory[501] = 3'b110;
        rom_memory[502] = 3'b110;
        rom_memory[503] = 3'b110;
        rom_memory[504] = 3'b110;
        rom_memory[505] = 3'b110;
        rom_memory[506] = 3'b110;
        rom_memory[507] = 3'b110;
        rom_memory[508] = 3'b110;
        rom_memory[509] = 3'b110;
        rom_memory[510] = 3'b110;
        rom_memory[511] = 3'b110;
        rom_memory[512] = 3'b110;
        rom_memory[513] = 3'b110;
        rom_memory[514] = 3'b110;
        rom_memory[515] = 3'b110;
        rom_memory[516] = 3'b110;
        rom_memory[517] = 3'b110;
        rom_memory[518] = 3'b110;
        rom_memory[519] = 3'b110;
        rom_memory[520] = 3'b110;
        rom_memory[521] = 3'b110;
        rom_memory[522] = 3'b110;
        rom_memory[523] = 3'b110;
        rom_memory[524] = 3'b110;
        rom_memory[525] = 3'b110;
        rom_memory[526] = 3'b110;
        rom_memory[527] = 3'b110;
        rom_memory[528] = 3'b110;
        rom_memory[529] = 3'b110;
        rom_memory[530] = 3'b110;
        rom_memory[531] = 3'b110;
        rom_memory[532] = 3'b110;
        rom_memory[533] = 3'b110;
        rom_memory[534] = 3'b110;
        rom_memory[535] = 3'b110;
        rom_memory[536] = 3'b110;
        rom_memory[537] = 3'b110;
        rom_memory[538] = 3'b110;
        rom_memory[539] = 3'b110;
        rom_memory[540] = 3'b110;
        rom_memory[541] = 3'b110;
        rom_memory[542] = 3'b110;
        rom_memory[543] = 3'b110;
        rom_memory[544] = 3'b110;
        rom_memory[545] = 3'b110;
        rom_memory[546] = 3'b110;
        rom_memory[547] = 3'b110;
        rom_memory[548] = 3'b110;
        rom_memory[549] = 3'b110;
        rom_memory[550] = 3'b110;
        rom_memory[551] = 3'b110;
        rom_memory[552] = 3'b110;
        rom_memory[553] = 3'b110;
        rom_memory[554] = 3'b110;
        rom_memory[555] = 3'b110;
        rom_memory[556] = 3'b110;
        rom_memory[557] = 3'b110;
        rom_memory[558] = 3'b110;
        rom_memory[559] = 3'b110;
        rom_memory[560] = 3'b110;
        rom_memory[561] = 3'b110;
        rom_memory[562] = 3'b110;
        rom_memory[563] = 3'b110;
        rom_memory[564] = 3'b110;
        rom_memory[565] = 3'b110;
        rom_memory[566] = 3'b110;
        rom_memory[567] = 3'b110;
        rom_memory[568] = 3'b110;
        rom_memory[569] = 3'b110;
        rom_memory[570] = 3'b110;
        rom_memory[571] = 3'b110;
        rom_memory[572] = 3'b110;
        rom_memory[573] = 3'b110;
        rom_memory[574] = 3'b110;
        rom_memory[575] = 3'b110;
        rom_memory[576] = 3'b110;
        rom_memory[577] = 3'b110;
        rom_memory[578] = 3'b110;
        rom_memory[579] = 3'b110;
        rom_memory[580] = 3'b110;
        rom_memory[581] = 3'b110;
        rom_memory[582] = 3'b110;
        rom_memory[583] = 3'b110;
        rom_memory[584] = 3'b110;
        rom_memory[585] = 3'b110;
        rom_memory[586] = 3'b110;
        rom_memory[587] = 3'b110;
        rom_memory[588] = 3'b110;
        rom_memory[589] = 3'b110;
        rom_memory[590] = 3'b110;
        rom_memory[591] = 3'b110;
        rom_memory[592] = 3'b110;
        rom_memory[593] = 3'b110;
        rom_memory[594] = 3'b110;
        rom_memory[595] = 3'b110;
        rom_memory[596] = 3'b110;
        rom_memory[597] = 3'b110;
        rom_memory[598] = 3'b110;
        rom_memory[599] = 3'b110;
        rom_memory[600] = 3'b110;
        rom_memory[601] = 3'b110;
        rom_memory[602] = 3'b110;
        rom_memory[603] = 3'b110;
        rom_memory[604] = 3'b110;
        rom_memory[605] = 3'b110;
        rom_memory[606] = 3'b110;
        rom_memory[607] = 3'b110;
        rom_memory[608] = 3'b110;
        rom_memory[609] = 3'b110;
        rom_memory[610] = 3'b110;
        rom_memory[611] = 3'b110;
        rom_memory[612] = 3'b110;
        rom_memory[613] = 3'b110;
        rom_memory[614] = 3'b110;
        rom_memory[615] = 3'b110;
        rom_memory[616] = 3'b110;
        rom_memory[617] = 3'b110;
        rom_memory[618] = 3'b110;
        rom_memory[619] = 3'b110;
        rom_memory[620] = 3'b110;
        rom_memory[621] = 3'b110;
        rom_memory[622] = 3'b110;
        rom_memory[623] = 3'b110;
        rom_memory[624] = 3'b110;
        rom_memory[625] = 3'b110;
        rom_memory[626] = 3'b110;
        rom_memory[627] = 3'b110;
        rom_memory[628] = 3'b110;
        rom_memory[629] = 3'b110;
        rom_memory[630] = 3'b110;
        rom_memory[631] = 3'b110;
        rom_memory[632] = 3'b110;
        rom_memory[633] = 3'b110;
        rom_memory[634] = 3'b110;
        rom_memory[635] = 3'b110;
        rom_memory[636] = 3'b110;
        rom_memory[637] = 3'b110;
        rom_memory[638] = 3'b100;
        rom_memory[639] = 3'b100;
        rom_memory[640] = 3'b100;
        rom_memory[641] = 3'b100;
        rom_memory[642] = 3'b100;
        rom_memory[643] = 3'b100;
        rom_memory[644] = 3'b100;
        rom_memory[645] = 3'b100;
        rom_memory[646] = 3'b100;
        rom_memory[647] = 3'b100;
        rom_memory[648] = 3'b100;
        rom_memory[649] = 3'b100;
        rom_memory[650] = 3'b100;
        rom_memory[651] = 3'b100;
        rom_memory[652] = 3'b100;
        rom_memory[653] = 3'b100;
        rom_memory[654] = 3'b100;
        rom_memory[655] = 3'b100;
        rom_memory[656] = 3'b100;
        rom_memory[657] = 3'b100;
        rom_memory[658] = 3'b100;
        rom_memory[659] = 3'b100;
        rom_memory[660] = 3'b100;
        rom_memory[661] = 3'b100;
        rom_memory[662] = 3'b100;
        rom_memory[663] = 3'b100;
        rom_memory[664] = 3'b100;
        rom_memory[665] = 3'b100;
        rom_memory[666] = 3'b100;
        rom_memory[667] = 3'b100;
        rom_memory[668] = 3'b100;
        rom_memory[669] = 3'b100;
        rom_memory[670] = 3'b100;
        rom_memory[671] = 3'b100;
        rom_memory[672] = 3'b100;
        rom_memory[673] = 3'b100;
        rom_memory[674] = 3'b100;
        rom_memory[675] = 3'b100;
        rom_memory[676] = 3'b100;
        rom_memory[677] = 3'b100;
        rom_memory[678] = 3'b100;
        rom_memory[679] = 3'b100;
        rom_memory[680] = 3'b100;
        rom_memory[681] = 3'b100;
        rom_memory[682] = 3'b100;
        rom_memory[683] = 3'b100;
        rom_memory[684] = 3'b100;
        rom_memory[685] = 3'b100;
        rom_memory[686] = 3'b100;
        rom_memory[687] = 3'b100;
        rom_memory[688] = 3'b100;
        rom_memory[689] = 3'b100;
        rom_memory[690] = 3'b100;
        rom_memory[691] = 3'b100;
        rom_memory[692] = 3'b100;
        rom_memory[693] = 3'b100;
        rom_memory[694] = 3'b100;
        rom_memory[695] = 3'b100;
        rom_memory[696] = 3'b100;
        rom_memory[697] = 3'b100;
        rom_memory[698] = 3'b100;
        rom_memory[699] = 3'b100;
        rom_memory[700] = 3'b100;
        rom_memory[701] = 3'b100;
        rom_memory[702] = 3'b100;
        rom_memory[703] = 3'b100;
        rom_memory[704] = 3'b100;
        rom_memory[705] = 3'b100;
        rom_memory[706] = 3'b100;
        rom_memory[707] = 3'b100;
        rom_memory[708] = 3'b100;
        rom_memory[709] = 3'b100;
        rom_memory[710] = 3'b100;
        rom_memory[711] = 3'b100;
        rom_memory[712] = 3'b100;
        rom_memory[713] = 3'b100;
        rom_memory[714] = 3'b100;
        rom_memory[715] = 3'b100;
        rom_memory[716] = 3'b100;
        rom_memory[717] = 3'b100;
        rom_memory[718] = 3'b100;
        rom_memory[719] = 3'b100;
        rom_memory[720] = 3'b110;
        rom_memory[721] = 3'b110;
        rom_memory[722] = 3'b110;
        rom_memory[723] = 3'b110;
        rom_memory[724] = 3'b110;
        rom_memory[725] = 3'b110;
        rom_memory[726] = 3'b110;
        rom_memory[727] = 3'b110;
        rom_memory[728] = 3'b110;
        rom_memory[729] = 3'b110;
        rom_memory[730] = 3'b110;
        rom_memory[731] = 3'b110;
        rom_memory[732] = 3'b110;
        rom_memory[733] = 3'b110;
        rom_memory[734] = 3'b110;
        rom_memory[735] = 3'b110;
        rom_memory[736] = 3'b110;
        rom_memory[737] = 3'b110;
        rom_memory[738] = 3'b110;
        rom_memory[739] = 3'b110;
        rom_memory[740] = 3'b110;
        rom_memory[741] = 3'b110;
        rom_memory[742] = 3'b110;
        rom_memory[743] = 3'b110;
        rom_memory[744] = 3'b110;
        rom_memory[745] = 3'b110;
        rom_memory[746] = 3'b110;
        rom_memory[747] = 3'b110;
        rom_memory[748] = 3'b110;
        rom_memory[749] = 3'b110;
        rom_memory[750] = 3'b110;
        rom_memory[751] = 3'b110;
        rom_memory[752] = 3'b110;
        rom_memory[753] = 3'b110;
        rom_memory[754] = 3'b110;
        rom_memory[755] = 3'b110;
        rom_memory[756] = 3'b110;
        rom_memory[757] = 3'b110;
        rom_memory[758] = 3'b110;
        rom_memory[759] = 3'b110;
        rom_memory[760] = 3'b110;
        rom_memory[761] = 3'b110;
        rom_memory[762] = 3'b110;
        rom_memory[763] = 3'b110;
        rom_memory[764] = 3'b110;
        rom_memory[765] = 3'b110;
        rom_memory[766] = 3'b110;
        rom_memory[767] = 3'b110;
        rom_memory[768] = 3'b110;
        rom_memory[769] = 3'b110;
        rom_memory[770] = 3'b110;
        rom_memory[771] = 3'b110;
        rom_memory[772] = 3'b110;
        rom_memory[773] = 3'b110;
        rom_memory[774] = 3'b110;
        rom_memory[775] = 3'b110;
        rom_memory[776] = 3'b110;
        rom_memory[777] = 3'b110;
        rom_memory[778] = 3'b110;
        rom_memory[779] = 3'b110;
        rom_memory[780] = 3'b110;
        rom_memory[781] = 3'b110;
        rom_memory[782] = 3'b110;
        rom_memory[783] = 3'b110;
        rom_memory[784] = 3'b110;
        rom_memory[785] = 3'b110;
        rom_memory[786] = 3'b110;
        rom_memory[787] = 3'b110;
        rom_memory[788] = 3'b110;
        rom_memory[789] = 3'b110;
        rom_memory[790] = 3'b110;
        rom_memory[791] = 3'b110;
        rom_memory[792] = 3'b110;
        rom_memory[793] = 3'b110;
        rom_memory[794] = 3'b110;
        rom_memory[795] = 3'b110;
        rom_memory[796] = 3'b110;
        rom_memory[797] = 3'b110;
        rom_memory[798] = 3'b110;
        rom_memory[799] = 3'b110;
        rom_memory[800] = 3'b110;
        rom_memory[801] = 3'b110;
        rom_memory[802] = 3'b110;
        rom_memory[803] = 3'b110;
        rom_memory[804] = 3'b110;
        rom_memory[805] = 3'b110;
        rom_memory[806] = 3'b110;
        rom_memory[807] = 3'b110;
        rom_memory[808] = 3'b110;
        rom_memory[809] = 3'b110;
        rom_memory[810] = 3'b110;
        rom_memory[811] = 3'b110;
        rom_memory[812] = 3'b110;
        rom_memory[813] = 3'b110;
        rom_memory[814] = 3'b110;
        rom_memory[815] = 3'b110;
        rom_memory[816] = 3'b110;
        rom_memory[817] = 3'b110;
        rom_memory[818] = 3'b110;
        rom_memory[819] = 3'b110;
        rom_memory[820] = 3'b110;
        rom_memory[821] = 3'b110;
        rom_memory[822] = 3'b110;
        rom_memory[823] = 3'b110;
        rom_memory[824] = 3'b110;
        rom_memory[825] = 3'b110;
        rom_memory[826] = 3'b110;
        rom_memory[827] = 3'b110;
        rom_memory[828] = 3'b110;
        rom_memory[829] = 3'b110;
        rom_memory[830] = 3'b110;
        rom_memory[831] = 3'b110;
        rom_memory[832] = 3'b110;
        rom_memory[833] = 3'b110;
        rom_memory[834] = 3'b110;
        rom_memory[835] = 3'b110;
        rom_memory[836] = 3'b110;
        rom_memory[837] = 3'b110;
        rom_memory[838] = 3'b110;
        rom_memory[839] = 3'b110;
        rom_memory[840] = 3'b110;
        rom_memory[841] = 3'b110;
        rom_memory[842] = 3'b110;
        rom_memory[843] = 3'b110;
        rom_memory[844] = 3'b110;
        rom_memory[845] = 3'b110;
        rom_memory[846] = 3'b110;
        rom_memory[847] = 3'b110;
        rom_memory[848] = 3'b110;
        rom_memory[849] = 3'b110;
        rom_memory[850] = 3'b110;
        rom_memory[851] = 3'b110;
        rom_memory[852] = 3'b110;
        rom_memory[853] = 3'b110;
        rom_memory[854] = 3'b110;
        rom_memory[855] = 3'b110;
        rom_memory[856] = 3'b110;
        rom_memory[857] = 3'b110;
        rom_memory[858] = 3'b110;
        rom_memory[859] = 3'b110;
        rom_memory[860] = 3'b110;
        rom_memory[861] = 3'b110;
        rom_memory[862] = 3'b110;
        rom_memory[863] = 3'b110;
        rom_memory[864] = 3'b110;
        rom_memory[865] = 3'b110;
        rom_memory[866] = 3'b110;
        rom_memory[867] = 3'b110;
        rom_memory[868] = 3'b110;
        rom_memory[869] = 3'b110;
        rom_memory[870] = 3'b110;
        rom_memory[871] = 3'b110;
        rom_memory[872] = 3'b110;
        rom_memory[873] = 3'b110;
        rom_memory[874] = 3'b110;
        rom_memory[875] = 3'b110;
        rom_memory[876] = 3'b110;
        rom_memory[877] = 3'b110;
        rom_memory[878] = 3'b110;
        rom_memory[879] = 3'b110;
        rom_memory[880] = 3'b100;
        rom_memory[881] = 3'b100;
        rom_memory[882] = 3'b100;
        rom_memory[883] = 3'b100;
        rom_memory[884] = 3'b100;
        rom_memory[885] = 3'b100;
        rom_memory[886] = 3'b100;
        rom_memory[887] = 3'b100;
        rom_memory[888] = 3'b100;
        rom_memory[889] = 3'b100;
        rom_memory[890] = 3'b100;
        rom_memory[891] = 3'b100;
        rom_memory[892] = 3'b100;
        rom_memory[893] = 3'b100;
        rom_memory[894] = 3'b100;
        rom_memory[895] = 3'b100;
        rom_memory[896] = 3'b100;
        rom_memory[897] = 3'b100;
        rom_memory[898] = 3'b100;
        rom_memory[899] = 3'b100;
        rom_memory[900] = 3'b100;
        rom_memory[901] = 3'b100;
        rom_memory[902] = 3'b100;
        rom_memory[903] = 3'b100;
        rom_memory[904] = 3'b100;
        rom_memory[905] = 3'b100;
        rom_memory[906] = 3'b100;
        rom_memory[907] = 3'b100;
        rom_memory[908] = 3'b100;
        rom_memory[909] = 3'b100;
        rom_memory[910] = 3'b100;
        rom_memory[911] = 3'b100;
        rom_memory[912] = 3'b100;
        rom_memory[913] = 3'b100;
        rom_memory[914] = 3'b100;
        rom_memory[915] = 3'b100;
        rom_memory[916] = 3'b100;
        rom_memory[917] = 3'b100;
        rom_memory[918] = 3'b100;
        rom_memory[919] = 3'b100;
        rom_memory[920] = 3'b100;
        rom_memory[921] = 3'b100;
        rom_memory[922] = 3'b100;
        rom_memory[923] = 3'b100;
        rom_memory[924] = 3'b100;
        rom_memory[925] = 3'b100;
        rom_memory[926] = 3'b100;
        rom_memory[927] = 3'b100;
        rom_memory[928] = 3'b100;
        rom_memory[929] = 3'b100;
        rom_memory[930] = 3'b100;
        rom_memory[931] = 3'b100;
        rom_memory[932] = 3'b100;
        rom_memory[933] = 3'b100;
        rom_memory[934] = 3'b100;
        rom_memory[935] = 3'b100;
        rom_memory[936] = 3'b100;
        rom_memory[937] = 3'b100;
        rom_memory[938] = 3'b100;
        rom_memory[939] = 3'b100;
        rom_memory[940] = 3'b100;
        rom_memory[941] = 3'b100;
        rom_memory[942] = 3'b100;
        rom_memory[943] = 3'b100;
        rom_memory[944] = 3'b100;
        rom_memory[945] = 3'b100;
        rom_memory[946] = 3'b100;
        rom_memory[947] = 3'b100;
        rom_memory[948] = 3'b100;
        rom_memory[949] = 3'b100;
        rom_memory[950] = 3'b100;
        rom_memory[951] = 3'b100;
        rom_memory[952] = 3'b100;
        rom_memory[953] = 3'b100;
        rom_memory[954] = 3'b100;
        rom_memory[955] = 3'b100;
        rom_memory[956] = 3'b100;
        rom_memory[957] = 3'b100;
        rom_memory[958] = 3'b100;
        rom_memory[959] = 3'b100;
        rom_memory[960] = 3'b110;
        rom_memory[961] = 3'b110;
        rom_memory[962] = 3'b110;
        rom_memory[963] = 3'b110;
        rom_memory[964] = 3'b110;
        rom_memory[965] = 3'b110;
        rom_memory[966] = 3'b110;
        rom_memory[967] = 3'b110;
        rom_memory[968] = 3'b110;
        rom_memory[969] = 3'b110;
        rom_memory[970] = 3'b110;
        rom_memory[971] = 3'b110;
        rom_memory[972] = 3'b110;
        rom_memory[973] = 3'b110;
        rom_memory[974] = 3'b110;
        rom_memory[975] = 3'b110;
        rom_memory[976] = 3'b110;
        rom_memory[977] = 3'b110;
        rom_memory[978] = 3'b110;
        rom_memory[979] = 3'b110;
        rom_memory[980] = 3'b110;
        rom_memory[981] = 3'b110;
        rom_memory[982] = 3'b110;
        rom_memory[983] = 3'b110;
        rom_memory[984] = 3'b110;
        rom_memory[985] = 3'b110;
        rom_memory[986] = 3'b110;
        rom_memory[987] = 3'b110;
        rom_memory[988] = 3'b110;
        rom_memory[989] = 3'b110;
        rom_memory[990] = 3'b110;
        rom_memory[991] = 3'b110;
        rom_memory[992] = 3'b110;
        rom_memory[993] = 3'b110;
        rom_memory[994] = 3'b110;
        rom_memory[995] = 3'b110;
        rom_memory[996] = 3'b110;
        rom_memory[997] = 3'b110;
        rom_memory[998] = 3'b110;
        rom_memory[999] = 3'b110;
        rom_memory[1000] = 3'b110;
        rom_memory[1001] = 3'b110;
        rom_memory[1002] = 3'b110;
        rom_memory[1003] = 3'b110;
        rom_memory[1004] = 3'b110;
        rom_memory[1005] = 3'b110;
        rom_memory[1006] = 3'b110;
        rom_memory[1007] = 3'b110;
        rom_memory[1008] = 3'b110;
        rom_memory[1009] = 3'b110;
        rom_memory[1010] = 3'b110;
        rom_memory[1011] = 3'b110;
        rom_memory[1012] = 3'b110;
        rom_memory[1013] = 3'b110;
        rom_memory[1014] = 3'b110;
        rom_memory[1015] = 3'b110;
        rom_memory[1016] = 3'b110;
        rom_memory[1017] = 3'b110;
        rom_memory[1018] = 3'b110;
        rom_memory[1019] = 3'b110;
        rom_memory[1020] = 3'b110;
        rom_memory[1021] = 3'b110;
        rom_memory[1022] = 3'b110;
        rom_memory[1023] = 3'b110;
        rom_memory[1024] = 3'b110;
        rom_memory[1025] = 3'b110;
        rom_memory[1026] = 3'b110;
        rom_memory[1027] = 3'b110;
        rom_memory[1028] = 3'b110;
        rom_memory[1029] = 3'b110;
        rom_memory[1030] = 3'b110;
        rom_memory[1031] = 3'b110;
        rom_memory[1032] = 3'b110;
        rom_memory[1033] = 3'b110;
        rom_memory[1034] = 3'b110;
        rom_memory[1035] = 3'b110;
        rom_memory[1036] = 3'b110;
        rom_memory[1037] = 3'b110;
        rom_memory[1038] = 3'b110;
        rom_memory[1039] = 3'b110;
        rom_memory[1040] = 3'b110;
        rom_memory[1041] = 3'b110;
        rom_memory[1042] = 3'b110;
        rom_memory[1043] = 3'b110;
        rom_memory[1044] = 3'b110;
        rom_memory[1045] = 3'b110;
        rom_memory[1046] = 3'b110;
        rom_memory[1047] = 3'b110;
        rom_memory[1048] = 3'b110;
        rom_memory[1049] = 3'b110;
        rom_memory[1050] = 3'b110;
        rom_memory[1051] = 3'b110;
        rom_memory[1052] = 3'b110;
        rom_memory[1053] = 3'b110;
        rom_memory[1054] = 3'b110;
        rom_memory[1055] = 3'b110;
        rom_memory[1056] = 3'b110;
        rom_memory[1057] = 3'b110;
        rom_memory[1058] = 3'b110;
        rom_memory[1059] = 3'b110;
        rom_memory[1060] = 3'b110;
        rom_memory[1061] = 3'b110;
        rom_memory[1062] = 3'b110;
        rom_memory[1063] = 3'b110;
        rom_memory[1064] = 3'b110;
        rom_memory[1065] = 3'b110;
        rom_memory[1066] = 3'b110;
        rom_memory[1067] = 3'b110;
        rom_memory[1068] = 3'b110;
        rom_memory[1069] = 3'b110;
        rom_memory[1070] = 3'b110;
        rom_memory[1071] = 3'b110;
        rom_memory[1072] = 3'b110;
        rom_memory[1073] = 3'b110;
        rom_memory[1074] = 3'b110;
        rom_memory[1075] = 3'b110;
        rom_memory[1076] = 3'b110;
        rom_memory[1077] = 3'b110;
        rom_memory[1078] = 3'b110;
        rom_memory[1079] = 3'b110;
        rom_memory[1080] = 3'b110;
        rom_memory[1081] = 3'b110;
        rom_memory[1082] = 3'b110;
        rom_memory[1083] = 3'b110;
        rom_memory[1084] = 3'b110;
        rom_memory[1085] = 3'b110;
        rom_memory[1086] = 3'b110;
        rom_memory[1087] = 3'b110;
        rom_memory[1088] = 3'b110;
        rom_memory[1089] = 3'b110;
        rom_memory[1090] = 3'b110;
        rom_memory[1091] = 3'b110;
        rom_memory[1092] = 3'b110;
        rom_memory[1093] = 3'b110;
        rom_memory[1094] = 3'b110;
        rom_memory[1095] = 3'b110;
        rom_memory[1096] = 3'b110;
        rom_memory[1097] = 3'b110;
        rom_memory[1098] = 3'b110;
        rom_memory[1099] = 3'b110;
        rom_memory[1100] = 3'b110;
        rom_memory[1101] = 3'b110;
        rom_memory[1102] = 3'b110;
        rom_memory[1103] = 3'b110;
        rom_memory[1104] = 3'b110;
        rom_memory[1105] = 3'b110;
        rom_memory[1106] = 3'b110;
        rom_memory[1107] = 3'b110;
        rom_memory[1108] = 3'b110;
        rom_memory[1109] = 3'b110;
        rom_memory[1110] = 3'b110;
        rom_memory[1111] = 3'b110;
        rom_memory[1112] = 3'b110;
        rom_memory[1113] = 3'b110;
        rom_memory[1114] = 3'b110;
        rom_memory[1115] = 3'b110;
        rom_memory[1116] = 3'b110;
        rom_memory[1117] = 3'b110;
        rom_memory[1118] = 3'b110;
        rom_memory[1119] = 3'b110;
        rom_memory[1120] = 3'b100;
        rom_memory[1121] = 3'b100;
        rom_memory[1122] = 3'b100;
        rom_memory[1123] = 3'b100;
        rom_memory[1124] = 3'b100;
        rom_memory[1125] = 3'b100;
        rom_memory[1126] = 3'b100;
        rom_memory[1127] = 3'b100;
        rom_memory[1128] = 3'b100;
        rom_memory[1129] = 3'b100;
        rom_memory[1130] = 3'b100;
        rom_memory[1131] = 3'b100;
        rom_memory[1132] = 3'b100;
        rom_memory[1133] = 3'b100;
        rom_memory[1134] = 3'b100;
        rom_memory[1135] = 3'b100;
        rom_memory[1136] = 3'b100;
        rom_memory[1137] = 3'b100;
        rom_memory[1138] = 3'b100;
        rom_memory[1139] = 3'b100;
        rom_memory[1140] = 3'b100;
        rom_memory[1141] = 3'b100;
        rom_memory[1142] = 3'b100;
        rom_memory[1143] = 3'b100;
        rom_memory[1144] = 3'b100;
        rom_memory[1145] = 3'b100;
        rom_memory[1146] = 3'b100;
        rom_memory[1147] = 3'b100;
        rom_memory[1148] = 3'b100;
        rom_memory[1149] = 3'b100;
        rom_memory[1150] = 3'b100;
        rom_memory[1151] = 3'b100;
        rom_memory[1152] = 3'b100;
        rom_memory[1153] = 3'b100;
        rom_memory[1154] = 3'b100;
        rom_memory[1155] = 3'b100;
        rom_memory[1156] = 3'b100;
        rom_memory[1157] = 3'b100;
        rom_memory[1158] = 3'b100;
        rom_memory[1159] = 3'b100;
        rom_memory[1160] = 3'b100;
        rom_memory[1161] = 3'b100;
        rom_memory[1162] = 3'b100;
        rom_memory[1163] = 3'b100;
        rom_memory[1164] = 3'b100;
        rom_memory[1165] = 3'b100;
        rom_memory[1166] = 3'b100;
        rom_memory[1167] = 3'b100;
        rom_memory[1168] = 3'b100;
        rom_memory[1169] = 3'b100;
        rom_memory[1170] = 3'b100;
        rom_memory[1171] = 3'b100;
        rom_memory[1172] = 3'b100;
        rom_memory[1173] = 3'b100;
        rom_memory[1174] = 3'b100;
        rom_memory[1175] = 3'b100;
        rom_memory[1176] = 3'b100;
        rom_memory[1177] = 3'b100;
        rom_memory[1178] = 3'b100;
        rom_memory[1179] = 3'b100;
        rom_memory[1180] = 3'b100;
        rom_memory[1181] = 3'b100;
        rom_memory[1182] = 3'b100;
        rom_memory[1183] = 3'b100;
        rom_memory[1184] = 3'b100;
        rom_memory[1185] = 3'b100;
        rom_memory[1186] = 3'b100;
        rom_memory[1187] = 3'b100;
        rom_memory[1188] = 3'b100;
        rom_memory[1189] = 3'b100;
        rom_memory[1190] = 3'b100;
        rom_memory[1191] = 3'b100;
        rom_memory[1192] = 3'b100;
        rom_memory[1193] = 3'b100;
        rom_memory[1194] = 3'b100;
        rom_memory[1195] = 3'b100;
        rom_memory[1196] = 3'b100;
        rom_memory[1197] = 3'b100;
        rom_memory[1198] = 3'b100;
        rom_memory[1199] = 3'b100;
        rom_memory[1200] = 3'b110;
        rom_memory[1201] = 3'b110;
        rom_memory[1202] = 3'b110;
        rom_memory[1203] = 3'b110;
        rom_memory[1204] = 3'b110;
        rom_memory[1205] = 3'b110;
        rom_memory[1206] = 3'b110;
        rom_memory[1207] = 3'b110;
        rom_memory[1208] = 3'b110;
        rom_memory[1209] = 3'b110;
        rom_memory[1210] = 3'b110;
        rom_memory[1211] = 3'b110;
        rom_memory[1212] = 3'b110;
        rom_memory[1213] = 3'b110;
        rom_memory[1214] = 3'b110;
        rom_memory[1215] = 3'b110;
        rom_memory[1216] = 3'b110;
        rom_memory[1217] = 3'b110;
        rom_memory[1218] = 3'b110;
        rom_memory[1219] = 3'b110;
        rom_memory[1220] = 3'b110;
        rom_memory[1221] = 3'b110;
        rom_memory[1222] = 3'b110;
        rom_memory[1223] = 3'b110;
        rom_memory[1224] = 3'b110;
        rom_memory[1225] = 3'b110;
        rom_memory[1226] = 3'b110;
        rom_memory[1227] = 3'b110;
        rom_memory[1228] = 3'b110;
        rom_memory[1229] = 3'b110;
        rom_memory[1230] = 3'b110;
        rom_memory[1231] = 3'b110;
        rom_memory[1232] = 3'b110;
        rom_memory[1233] = 3'b110;
        rom_memory[1234] = 3'b110;
        rom_memory[1235] = 3'b110;
        rom_memory[1236] = 3'b110;
        rom_memory[1237] = 3'b110;
        rom_memory[1238] = 3'b110;
        rom_memory[1239] = 3'b110;
        rom_memory[1240] = 3'b110;
        rom_memory[1241] = 3'b110;
        rom_memory[1242] = 3'b110;
        rom_memory[1243] = 3'b110;
        rom_memory[1244] = 3'b110;
        rom_memory[1245] = 3'b110;
        rom_memory[1246] = 3'b110;
        rom_memory[1247] = 3'b110;
        rom_memory[1248] = 3'b110;
        rom_memory[1249] = 3'b110;
        rom_memory[1250] = 3'b110;
        rom_memory[1251] = 3'b110;
        rom_memory[1252] = 3'b110;
        rom_memory[1253] = 3'b110;
        rom_memory[1254] = 3'b110;
        rom_memory[1255] = 3'b110;
        rom_memory[1256] = 3'b110;
        rom_memory[1257] = 3'b110;
        rom_memory[1258] = 3'b110;
        rom_memory[1259] = 3'b110;
        rom_memory[1260] = 3'b110;
        rom_memory[1261] = 3'b110;
        rom_memory[1262] = 3'b110;
        rom_memory[1263] = 3'b110;
        rom_memory[1264] = 3'b110;
        rom_memory[1265] = 3'b110;
        rom_memory[1266] = 3'b110;
        rom_memory[1267] = 3'b110;
        rom_memory[1268] = 3'b110;
        rom_memory[1269] = 3'b110;
        rom_memory[1270] = 3'b110;
        rom_memory[1271] = 3'b110;
        rom_memory[1272] = 3'b110;
        rom_memory[1273] = 3'b110;
        rom_memory[1274] = 3'b110;
        rom_memory[1275] = 3'b110;
        rom_memory[1276] = 3'b110;
        rom_memory[1277] = 3'b110;
        rom_memory[1278] = 3'b110;
        rom_memory[1279] = 3'b110;
        rom_memory[1280] = 3'b110;
        rom_memory[1281] = 3'b110;
        rom_memory[1282] = 3'b110;
        rom_memory[1283] = 3'b110;
        rom_memory[1284] = 3'b110;
        rom_memory[1285] = 3'b110;
        rom_memory[1286] = 3'b110;
        rom_memory[1287] = 3'b110;
        rom_memory[1288] = 3'b110;
        rom_memory[1289] = 3'b110;
        rom_memory[1290] = 3'b110;
        rom_memory[1291] = 3'b110;
        rom_memory[1292] = 3'b110;
        rom_memory[1293] = 3'b110;
        rom_memory[1294] = 3'b110;
        rom_memory[1295] = 3'b110;
        rom_memory[1296] = 3'b110;
        rom_memory[1297] = 3'b110;
        rom_memory[1298] = 3'b110;
        rom_memory[1299] = 3'b110;
        rom_memory[1300] = 3'b110;
        rom_memory[1301] = 3'b110;
        rom_memory[1302] = 3'b110;
        rom_memory[1303] = 3'b110;
        rom_memory[1304] = 3'b110;
        rom_memory[1305] = 3'b110;
        rom_memory[1306] = 3'b110;
        rom_memory[1307] = 3'b110;
        rom_memory[1308] = 3'b110;
        rom_memory[1309] = 3'b110;
        rom_memory[1310] = 3'b110;
        rom_memory[1311] = 3'b110;
        rom_memory[1312] = 3'b110;
        rom_memory[1313] = 3'b110;
        rom_memory[1314] = 3'b110;
        rom_memory[1315] = 3'b110;
        rom_memory[1316] = 3'b110;
        rom_memory[1317] = 3'b110;
        rom_memory[1318] = 3'b110;
        rom_memory[1319] = 3'b110;
        rom_memory[1320] = 3'b110;
        rom_memory[1321] = 3'b110;
        rom_memory[1322] = 3'b110;
        rom_memory[1323] = 3'b110;
        rom_memory[1324] = 3'b110;
        rom_memory[1325] = 3'b110;
        rom_memory[1326] = 3'b110;
        rom_memory[1327] = 3'b110;
        rom_memory[1328] = 3'b110;
        rom_memory[1329] = 3'b110;
        rom_memory[1330] = 3'b110;
        rom_memory[1331] = 3'b110;
        rom_memory[1332] = 3'b110;
        rom_memory[1333] = 3'b110;
        rom_memory[1334] = 3'b110;
        rom_memory[1335] = 3'b110;
        rom_memory[1336] = 3'b110;
        rom_memory[1337] = 3'b110;
        rom_memory[1338] = 3'b110;
        rom_memory[1339] = 3'b110;
        rom_memory[1340] = 3'b110;
        rom_memory[1341] = 3'b110;
        rom_memory[1342] = 3'b110;
        rom_memory[1343] = 3'b110;
        rom_memory[1344] = 3'b110;
        rom_memory[1345] = 3'b110;
        rom_memory[1346] = 3'b110;
        rom_memory[1347] = 3'b110;
        rom_memory[1348] = 3'b110;
        rom_memory[1349] = 3'b110;
        rom_memory[1350] = 3'b110;
        rom_memory[1351] = 3'b110;
        rom_memory[1352] = 3'b110;
        rom_memory[1353] = 3'b110;
        rom_memory[1354] = 3'b110;
        rom_memory[1355] = 3'b110;
        rom_memory[1356] = 3'b110;
        rom_memory[1357] = 3'b110;
        rom_memory[1358] = 3'b110;
        rom_memory[1359] = 3'b110;
        rom_memory[1360] = 3'b100;
        rom_memory[1361] = 3'b100;
        rom_memory[1362] = 3'b100;
        rom_memory[1363] = 3'b100;
        rom_memory[1364] = 3'b100;
        rom_memory[1365] = 3'b100;
        rom_memory[1366] = 3'b100;
        rom_memory[1367] = 3'b100;
        rom_memory[1368] = 3'b100;
        rom_memory[1369] = 3'b100;
        rom_memory[1370] = 3'b100;
        rom_memory[1371] = 3'b100;
        rom_memory[1372] = 3'b100;
        rom_memory[1373] = 3'b100;
        rom_memory[1374] = 3'b100;
        rom_memory[1375] = 3'b100;
        rom_memory[1376] = 3'b100;
        rom_memory[1377] = 3'b100;
        rom_memory[1378] = 3'b100;
        rom_memory[1379] = 3'b100;
        rom_memory[1380] = 3'b100;
        rom_memory[1381] = 3'b100;
        rom_memory[1382] = 3'b100;
        rom_memory[1383] = 3'b100;
        rom_memory[1384] = 3'b100;
        rom_memory[1385] = 3'b100;
        rom_memory[1386] = 3'b100;
        rom_memory[1387] = 3'b100;
        rom_memory[1388] = 3'b100;
        rom_memory[1389] = 3'b100;
        rom_memory[1390] = 3'b100;
        rom_memory[1391] = 3'b100;
        rom_memory[1392] = 3'b100;
        rom_memory[1393] = 3'b100;
        rom_memory[1394] = 3'b100;
        rom_memory[1395] = 3'b100;
        rom_memory[1396] = 3'b100;
        rom_memory[1397] = 3'b100;
        rom_memory[1398] = 3'b100;
        rom_memory[1399] = 3'b100;
        rom_memory[1400] = 3'b100;
        rom_memory[1401] = 3'b100;
        rom_memory[1402] = 3'b100;
        rom_memory[1403] = 3'b100;
        rom_memory[1404] = 3'b100;
        rom_memory[1405] = 3'b100;
        rom_memory[1406] = 3'b100;
        rom_memory[1407] = 3'b100;
        rom_memory[1408] = 3'b100;
        rom_memory[1409] = 3'b100;
        rom_memory[1410] = 3'b100;
        rom_memory[1411] = 3'b100;
        rom_memory[1412] = 3'b100;
        rom_memory[1413] = 3'b100;
        rom_memory[1414] = 3'b100;
        rom_memory[1415] = 3'b100;
        rom_memory[1416] = 3'b100;
        rom_memory[1417] = 3'b100;
        rom_memory[1418] = 3'b100;
        rom_memory[1419] = 3'b100;
        rom_memory[1420] = 3'b100;
        rom_memory[1421] = 3'b100;
        rom_memory[1422] = 3'b100;
        rom_memory[1423] = 3'b100;
        rom_memory[1424] = 3'b100;
        rom_memory[1425] = 3'b100;
        rom_memory[1426] = 3'b100;
        rom_memory[1427] = 3'b100;
        rom_memory[1428] = 3'b100;
        rom_memory[1429] = 3'b100;
        rom_memory[1430] = 3'b100;
        rom_memory[1431] = 3'b100;
        rom_memory[1432] = 3'b100;
        rom_memory[1433] = 3'b100;
        rom_memory[1434] = 3'b100;
        rom_memory[1435] = 3'b100;
        rom_memory[1436] = 3'b100;
        rom_memory[1437] = 3'b100;
        rom_memory[1438] = 3'b100;
        rom_memory[1439] = 3'b100;
        rom_memory[1440] = 3'b110;
        rom_memory[1441] = 3'b110;
        rom_memory[1442] = 3'b110;
        rom_memory[1443] = 3'b110;
        rom_memory[1444] = 3'b110;
        rom_memory[1445] = 3'b110;
        rom_memory[1446] = 3'b110;
        rom_memory[1447] = 3'b110;
        rom_memory[1448] = 3'b110;
        rom_memory[1449] = 3'b110;
        rom_memory[1450] = 3'b110;
        rom_memory[1451] = 3'b110;
        rom_memory[1452] = 3'b110;
        rom_memory[1453] = 3'b110;
        rom_memory[1454] = 3'b110;
        rom_memory[1455] = 3'b110;
        rom_memory[1456] = 3'b110;
        rom_memory[1457] = 3'b110;
        rom_memory[1458] = 3'b110;
        rom_memory[1459] = 3'b110;
        rom_memory[1460] = 3'b110;
        rom_memory[1461] = 3'b110;
        rom_memory[1462] = 3'b110;
        rom_memory[1463] = 3'b110;
        rom_memory[1464] = 3'b110;
        rom_memory[1465] = 3'b110;
        rom_memory[1466] = 3'b110;
        rom_memory[1467] = 3'b110;
        rom_memory[1468] = 3'b110;
        rom_memory[1469] = 3'b110;
        rom_memory[1470] = 3'b110;
        rom_memory[1471] = 3'b110;
        rom_memory[1472] = 3'b110;
        rom_memory[1473] = 3'b110;
        rom_memory[1474] = 3'b110;
        rom_memory[1475] = 3'b110;
        rom_memory[1476] = 3'b110;
        rom_memory[1477] = 3'b110;
        rom_memory[1478] = 3'b110;
        rom_memory[1479] = 3'b110;
        rom_memory[1480] = 3'b110;
        rom_memory[1481] = 3'b110;
        rom_memory[1482] = 3'b110;
        rom_memory[1483] = 3'b110;
        rom_memory[1484] = 3'b110;
        rom_memory[1485] = 3'b110;
        rom_memory[1486] = 3'b110;
        rom_memory[1487] = 3'b110;
        rom_memory[1488] = 3'b110;
        rom_memory[1489] = 3'b110;
        rom_memory[1490] = 3'b110;
        rom_memory[1491] = 3'b110;
        rom_memory[1492] = 3'b110;
        rom_memory[1493] = 3'b110;
        rom_memory[1494] = 3'b110;
        rom_memory[1495] = 3'b110;
        rom_memory[1496] = 3'b110;
        rom_memory[1497] = 3'b110;
        rom_memory[1498] = 3'b110;
        rom_memory[1499] = 3'b110;
        rom_memory[1500] = 3'b110;
        rom_memory[1501] = 3'b110;
        rom_memory[1502] = 3'b110;
        rom_memory[1503] = 3'b110;
        rom_memory[1504] = 3'b110;
        rom_memory[1505] = 3'b110;
        rom_memory[1506] = 3'b110;
        rom_memory[1507] = 3'b110;
        rom_memory[1508] = 3'b110;
        rom_memory[1509] = 3'b110;
        rom_memory[1510] = 3'b110;
        rom_memory[1511] = 3'b110;
        rom_memory[1512] = 3'b110;
        rom_memory[1513] = 3'b110;
        rom_memory[1514] = 3'b110;
        rom_memory[1515] = 3'b110;
        rom_memory[1516] = 3'b110;
        rom_memory[1517] = 3'b110;
        rom_memory[1518] = 3'b110;
        rom_memory[1519] = 3'b110;
        rom_memory[1520] = 3'b110;
        rom_memory[1521] = 3'b110;
        rom_memory[1522] = 3'b110;
        rom_memory[1523] = 3'b110;
        rom_memory[1524] = 3'b110;
        rom_memory[1525] = 3'b110;
        rom_memory[1526] = 3'b110;
        rom_memory[1527] = 3'b110;
        rom_memory[1528] = 3'b110;
        rom_memory[1529] = 3'b110;
        rom_memory[1530] = 3'b110;
        rom_memory[1531] = 3'b110;
        rom_memory[1532] = 3'b110;
        rom_memory[1533] = 3'b110;
        rom_memory[1534] = 3'b110;
        rom_memory[1535] = 3'b110;
        rom_memory[1536] = 3'b110;
        rom_memory[1537] = 3'b110;
        rom_memory[1538] = 3'b110;
        rom_memory[1539] = 3'b110;
        rom_memory[1540] = 3'b110;
        rom_memory[1541] = 3'b110;
        rom_memory[1542] = 3'b110;
        rom_memory[1543] = 3'b110;
        rom_memory[1544] = 3'b110;
        rom_memory[1545] = 3'b110;
        rom_memory[1546] = 3'b110;
        rom_memory[1547] = 3'b110;
        rom_memory[1548] = 3'b110;
        rom_memory[1549] = 3'b110;
        rom_memory[1550] = 3'b110;
        rom_memory[1551] = 3'b110;
        rom_memory[1552] = 3'b110;
        rom_memory[1553] = 3'b110;
        rom_memory[1554] = 3'b110;
        rom_memory[1555] = 3'b110;
        rom_memory[1556] = 3'b110;
        rom_memory[1557] = 3'b110;
        rom_memory[1558] = 3'b110;
        rom_memory[1559] = 3'b110;
        rom_memory[1560] = 3'b110;
        rom_memory[1561] = 3'b110;
        rom_memory[1562] = 3'b110;
        rom_memory[1563] = 3'b110;
        rom_memory[1564] = 3'b110;
        rom_memory[1565] = 3'b110;
        rom_memory[1566] = 3'b110;
        rom_memory[1567] = 3'b110;
        rom_memory[1568] = 3'b110;
        rom_memory[1569] = 3'b110;
        rom_memory[1570] = 3'b110;
        rom_memory[1571] = 3'b110;
        rom_memory[1572] = 3'b110;
        rom_memory[1573] = 3'b110;
        rom_memory[1574] = 3'b110;
        rom_memory[1575] = 3'b110;
        rom_memory[1576] = 3'b110;
        rom_memory[1577] = 3'b110;
        rom_memory[1578] = 3'b110;
        rom_memory[1579] = 3'b110;
        rom_memory[1580] = 3'b110;
        rom_memory[1581] = 3'b110;
        rom_memory[1582] = 3'b110;
        rom_memory[1583] = 3'b110;
        rom_memory[1584] = 3'b110;
        rom_memory[1585] = 3'b110;
        rom_memory[1586] = 3'b110;
        rom_memory[1587] = 3'b110;
        rom_memory[1588] = 3'b110;
        rom_memory[1589] = 3'b110;
        rom_memory[1590] = 3'b110;
        rom_memory[1591] = 3'b110;
        rom_memory[1592] = 3'b110;
        rom_memory[1593] = 3'b110;
        rom_memory[1594] = 3'b110;
        rom_memory[1595] = 3'b110;
        rom_memory[1596] = 3'b110;
        rom_memory[1597] = 3'b110;
        rom_memory[1598] = 3'b110;
        rom_memory[1599] = 3'b110;
        rom_memory[1600] = 3'b110;
        rom_memory[1601] = 3'b100;
        rom_memory[1602] = 3'b100;
        rom_memory[1603] = 3'b100;
        rom_memory[1604] = 3'b100;
        rom_memory[1605] = 3'b100;
        rom_memory[1606] = 3'b100;
        rom_memory[1607] = 3'b100;
        rom_memory[1608] = 3'b100;
        rom_memory[1609] = 3'b100;
        rom_memory[1610] = 3'b100;
        rom_memory[1611] = 3'b100;
        rom_memory[1612] = 3'b100;
        rom_memory[1613] = 3'b100;
        rom_memory[1614] = 3'b100;
        rom_memory[1615] = 3'b100;
        rom_memory[1616] = 3'b100;
        rom_memory[1617] = 3'b100;
        rom_memory[1618] = 3'b100;
        rom_memory[1619] = 3'b100;
        rom_memory[1620] = 3'b100;
        rom_memory[1621] = 3'b100;
        rom_memory[1622] = 3'b100;
        rom_memory[1623] = 3'b100;
        rom_memory[1624] = 3'b100;
        rom_memory[1625] = 3'b100;
        rom_memory[1626] = 3'b100;
        rom_memory[1627] = 3'b100;
        rom_memory[1628] = 3'b100;
        rom_memory[1629] = 3'b100;
        rom_memory[1630] = 3'b100;
        rom_memory[1631] = 3'b100;
        rom_memory[1632] = 3'b100;
        rom_memory[1633] = 3'b100;
        rom_memory[1634] = 3'b100;
        rom_memory[1635] = 3'b100;
        rom_memory[1636] = 3'b100;
        rom_memory[1637] = 3'b100;
        rom_memory[1638] = 3'b100;
        rom_memory[1639] = 3'b100;
        rom_memory[1640] = 3'b100;
        rom_memory[1641] = 3'b100;
        rom_memory[1642] = 3'b100;
        rom_memory[1643] = 3'b100;
        rom_memory[1644] = 3'b100;
        rom_memory[1645] = 3'b100;
        rom_memory[1646] = 3'b100;
        rom_memory[1647] = 3'b100;
        rom_memory[1648] = 3'b100;
        rom_memory[1649] = 3'b100;
        rom_memory[1650] = 3'b100;
        rom_memory[1651] = 3'b100;
        rom_memory[1652] = 3'b100;
        rom_memory[1653] = 3'b100;
        rom_memory[1654] = 3'b100;
        rom_memory[1655] = 3'b100;
        rom_memory[1656] = 3'b100;
        rom_memory[1657] = 3'b100;
        rom_memory[1658] = 3'b100;
        rom_memory[1659] = 3'b100;
        rom_memory[1660] = 3'b100;
        rom_memory[1661] = 3'b100;
        rom_memory[1662] = 3'b100;
        rom_memory[1663] = 3'b100;
        rom_memory[1664] = 3'b100;
        rom_memory[1665] = 3'b100;
        rom_memory[1666] = 3'b100;
        rom_memory[1667] = 3'b100;
        rom_memory[1668] = 3'b100;
        rom_memory[1669] = 3'b100;
        rom_memory[1670] = 3'b100;
        rom_memory[1671] = 3'b100;
        rom_memory[1672] = 3'b100;
        rom_memory[1673] = 3'b100;
        rom_memory[1674] = 3'b100;
        rom_memory[1675] = 3'b100;
        rom_memory[1676] = 3'b100;
        rom_memory[1677] = 3'b100;
        rom_memory[1678] = 3'b100;
        rom_memory[1679] = 3'b100;
        rom_memory[1680] = 3'b110;
        rom_memory[1681] = 3'b110;
        rom_memory[1682] = 3'b110;
        rom_memory[1683] = 3'b110;
        rom_memory[1684] = 3'b110;
        rom_memory[1685] = 3'b110;
        rom_memory[1686] = 3'b110;
        rom_memory[1687] = 3'b110;
        rom_memory[1688] = 3'b110;
        rom_memory[1689] = 3'b110;
        rom_memory[1690] = 3'b110;
        rom_memory[1691] = 3'b110;
        rom_memory[1692] = 3'b110;
        rom_memory[1693] = 3'b110;
        rom_memory[1694] = 3'b110;
        rom_memory[1695] = 3'b110;
        rom_memory[1696] = 3'b110;
        rom_memory[1697] = 3'b110;
        rom_memory[1698] = 3'b110;
        rom_memory[1699] = 3'b110;
        rom_memory[1700] = 3'b110;
        rom_memory[1701] = 3'b110;
        rom_memory[1702] = 3'b110;
        rom_memory[1703] = 3'b110;
        rom_memory[1704] = 3'b110;
        rom_memory[1705] = 3'b110;
        rom_memory[1706] = 3'b110;
        rom_memory[1707] = 3'b110;
        rom_memory[1708] = 3'b110;
        rom_memory[1709] = 3'b110;
        rom_memory[1710] = 3'b110;
        rom_memory[1711] = 3'b110;
        rom_memory[1712] = 3'b110;
        rom_memory[1713] = 3'b110;
        rom_memory[1714] = 3'b110;
        rom_memory[1715] = 3'b110;
        rom_memory[1716] = 3'b110;
        rom_memory[1717] = 3'b110;
        rom_memory[1718] = 3'b110;
        rom_memory[1719] = 3'b110;
        rom_memory[1720] = 3'b110;
        rom_memory[1721] = 3'b110;
        rom_memory[1722] = 3'b110;
        rom_memory[1723] = 3'b110;
        rom_memory[1724] = 3'b110;
        rom_memory[1725] = 3'b110;
        rom_memory[1726] = 3'b110;
        rom_memory[1727] = 3'b110;
        rom_memory[1728] = 3'b110;
        rom_memory[1729] = 3'b110;
        rom_memory[1730] = 3'b110;
        rom_memory[1731] = 3'b110;
        rom_memory[1732] = 3'b110;
        rom_memory[1733] = 3'b110;
        rom_memory[1734] = 3'b110;
        rom_memory[1735] = 3'b110;
        rom_memory[1736] = 3'b110;
        rom_memory[1737] = 3'b110;
        rom_memory[1738] = 3'b110;
        rom_memory[1739] = 3'b110;
        rom_memory[1740] = 3'b110;
        rom_memory[1741] = 3'b110;
        rom_memory[1742] = 3'b110;
        rom_memory[1743] = 3'b110;
        rom_memory[1744] = 3'b110;
        rom_memory[1745] = 3'b110;
        rom_memory[1746] = 3'b110;
        rom_memory[1747] = 3'b110;
        rom_memory[1748] = 3'b110;
        rom_memory[1749] = 3'b110;
        rom_memory[1750] = 3'b110;
        rom_memory[1751] = 3'b110;
        rom_memory[1752] = 3'b110;
        rom_memory[1753] = 3'b110;
        rom_memory[1754] = 3'b110;
        rom_memory[1755] = 3'b110;
        rom_memory[1756] = 3'b110;
        rom_memory[1757] = 3'b110;
        rom_memory[1758] = 3'b110;
        rom_memory[1759] = 3'b110;
        rom_memory[1760] = 3'b110;
        rom_memory[1761] = 3'b110;
        rom_memory[1762] = 3'b110;
        rom_memory[1763] = 3'b110;
        rom_memory[1764] = 3'b110;
        rom_memory[1765] = 3'b110;
        rom_memory[1766] = 3'b110;
        rom_memory[1767] = 3'b110;
        rom_memory[1768] = 3'b110;
        rom_memory[1769] = 3'b110;
        rom_memory[1770] = 3'b110;
        rom_memory[1771] = 3'b110;
        rom_memory[1772] = 3'b110;
        rom_memory[1773] = 3'b110;
        rom_memory[1774] = 3'b110;
        rom_memory[1775] = 3'b110;
        rom_memory[1776] = 3'b110;
        rom_memory[1777] = 3'b110;
        rom_memory[1778] = 3'b110;
        rom_memory[1779] = 3'b110;
        rom_memory[1780] = 3'b110;
        rom_memory[1781] = 3'b110;
        rom_memory[1782] = 3'b110;
        rom_memory[1783] = 3'b110;
        rom_memory[1784] = 3'b110;
        rom_memory[1785] = 3'b110;
        rom_memory[1786] = 3'b110;
        rom_memory[1787] = 3'b110;
        rom_memory[1788] = 3'b110;
        rom_memory[1789] = 3'b110;
        rom_memory[1790] = 3'b110;
        rom_memory[1791] = 3'b110;
        rom_memory[1792] = 3'b110;
        rom_memory[1793] = 3'b110;
        rom_memory[1794] = 3'b110;
        rom_memory[1795] = 3'b110;
        rom_memory[1796] = 3'b110;
        rom_memory[1797] = 3'b110;
        rom_memory[1798] = 3'b110;
        rom_memory[1799] = 3'b110;
        rom_memory[1800] = 3'b110;
        rom_memory[1801] = 3'b110;
        rom_memory[1802] = 3'b110;
        rom_memory[1803] = 3'b110;
        rom_memory[1804] = 3'b110;
        rom_memory[1805] = 3'b110;
        rom_memory[1806] = 3'b110;
        rom_memory[1807] = 3'b110;
        rom_memory[1808] = 3'b110;
        rom_memory[1809] = 3'b110;
        rom_memory[1810] = 3'b110;
        rom_memory[1811] = 3'b110;
        rom_memory[1812] = 3'b110;
        rom_memory[1813] = 3'b110;
        rom_memory[1814] = 3'b110;
        rom_memory[1815] = 3'b110;
        rom_memory[1816] = 3'b110;
        rom_memory[1817] = 3'b110;
        rom_memory[1818] = 3'b110;
        rom_memory[1819] = 3'b110;
        rom_memory[1820] = 3'b110;
        rom_memory[1821] = 3'b110;
        rom_memory[1822] = 3'b110;
        rom_memory[1823] = 3'b110;
        rom_memory[1824] = 3'b110;
        rom_memory[1825] = 3'b110;
        rom_memory[1826] = 3'b110;
        rom_memory[1827] = 3'b110;
        rom_memory[1828] = 3'b110;
        rom_memory[1829] = 3'b110;
        rom_memory[1830] = 3'b110;
        rom_memory[1831] = 3'b110;
        rom_memory[1832] = 3'b110;
        rom_memory[1833] = 3'b110;
        rom_memory[1834] = 3'b110;
        rom_memory[1835] = 3'b110;
        rom_memory[1836] = 3'b110;
        rom_memory[1837] = 3'b110;
        rom_memory[1838] = 3'b110;
        rom_memory[1839] = 3'b110;
        rom_memory[1840] = 3'b110;
        rom_memory[1841] = 3'b100;
        rom_memory[1842] = 3'b100;
        rom_memory[1843] = 3'b100;
        rom_memory[1844] = 3'b100;
        rom_memory[1845] = 3'b100;
        rom_memory[1846] = 3'b100;
        rom_memory[1847] = 3'b100;
        rom_memory[1848] = 3'b100;
        rom_memory[1849] = 3'b100;
        rom_memory[1850] = 3'b100;
        rom_memory[1851] = 3'b100;
        rom_memory[1852] = 3'b100;
        rom_memory[1853] = 3'b100;
        rom_memory[1854] = 3'b100;
        rom_memory[1855] = 3'b100;
        rom_memory[1856] = 3'b100;
        rom_memory[1857] = 3'b100;
        rom_memory[1858] = 3'b100;
        rom_memory[1859] = 3'b100;
        rom_memory[1860] = 3'b100;
        rom_memory[1861] = 3'b100;
        rom_memory[1862] = 3'b100;
        rom_memory[1863] = 3'b100;
        rom_memory[1864] = 3'b100;
        rom_memory[1865] = 3'b100;
        rom_memory[1866] = 3'b100;
        rom_memory[1867] = 3'b100;
        rom_memory[1868] = 3'b100;
        rom_memory[1869] = 3'b100;
        rom_memory[1870] = 3'b100;
        rom_memory[1871] = 3'b100;
        rom_memory[1872] = 3'b100;
        rom_memory[1873] = 3'b100;
        rom_memory[1874] = 3'b100;
        rom_memory[1875] = 3'b100;
        rom_memory[1876] = 3'b100;
        rom_memory[1877] = 3'b100;
        rom_memory[1878] = 3'b100;
        rom_memory[1879] = 3'b100;
        rom_memory[1880] = 3'b100;
        rom_memory[1881] = 3'b100;
        rom_memory[1882] = 3'b100;
        rom_memory[1883] = 3'b100;
        rom_memory[1884] = 3'b100;
        rom_memory[1885] = 3'b100;
        rom_memory[1886] = 3'b100;
        rom_memory[1887] = 3'b100;
        rom_memory[1888] = 3'b100;
        rom_memory[1889] = 3'b100;
        rom_memory[1890] = 3'b100;
        rom_memory[1891] = 3'b100;
        rom_memory[1892] = 3'b100;
        rom_memory[1893] = 3'b100;
        rom_memory[1894] = 3'b100;
        rom_memory[1895] = 3'b100;
        rom_memory[1896] = 3'b100;
        rom_memory[1897] = 3'b100;
        rom_memory[1898] = 3'b100;
        rom_memory[1899] = 3'b100;
        rom_memory[1900] = 3'b100;
        rom_memory[1901] = 3'b100;
        rom_memory[1902] = 3'b100;
        rom_memory[1903] = 3'b100;
        rom_memory[1904] = 3'b100;
        rom_memory[1905] = 3'b100;
        rom_memory[1906] = 3'b100;
        rom_memory[1907] = 3'b100;
        rom_memory[1908] = 3'b100;
        rom_memory[1909] = 3'b100;
        rom_memory[1910] = 3'b100;
        rom_memory[1911] = 3'b100;
        rom_memory[1912] = 3'b100;
        rom_memory[1913] = 3'b100;
        rom_memory[1914] = 3'b100;
        rom_memory[1915] = 3'b100;
        rom_memory[1916] = 3'b100;
        rom_memory[1917] = 3'b100;
        rom_memory[1918] = 3'b100;
        rom_memory[1919] = 3'b100;
        rom_memory[1920] = 3'b110;
        rom_memory[1921] = 3'b110;
        rom_memory[1922] = 3'b110;
        rom_memory[1923] = 3'b110;
        rom_memory[1924] = 3'b110;
        rom_memory[1925] = 3'b110;
        rom_memory[1926] = 3'b110;
        rom_memory[1927] = 3'b110;
        rom_memory[1928] = 3'b110;
        rom_memory[1929] = 3'b110;
        rom_memory[1930] = 3'b110;
        rom_memory[1931] = 3'b110;
        rom_memory[1932] = 3'b110;
        rom_memory[1933] = 3'b110;
        rom_memory[1934] = 3'b110;
        rom_memory[1935] = 3'b110;
        rom_memory[1936] = 3'b110;
        rom_memory[1937] = 3'b110;
        rom_memory[1938] = 3'b110;
        rom_memory[1939] = 3'b110;
        rom_memory[1940] = 3'b110;
        rom_memory[1941] = 3'b110;
        rom_memory[1942] = 3'b110;
        rom_memory[1943] = 3'b110;
        rom_memory[1944] = 3'b110;
        rom_memory[1945] = 3'b110;
        rom_memory[1946] = 3'b110;
        rom_memory[1947] = 3'b110;
        rom_memory[1948] = 3'b110;
        rom_memory[1949] = 3'b110;
        rom_memory[1950] = 3'b110;
        rom_memory[1951] = 3'b110;
        rom_memory[1952] = 3'b110;
        rom_memory[1953] = 3'b110;
        rom_memory[1954] = 3'b110;
        rom_memory[1955] = 3'b110;
        rom_memory[1956] = 3'b110;
        rom_memory[1957] = 3'b110;
        rom_memory[1958] = 3'b110;
        rom_memory[1959] = 3'b110;
        rom_memory[1960] = 3'b110;
        rom_memory[1961] = 3'b110;
        rom_memory[1962] = 3'b110;
        rom_memory[1963] = 3'b110;
        rom_memory[1964] = 3'b110;
        rom_memory[1965] = 3'b110;
        rom_memory[1966] = 3'b110;
        rom_memory[1967] = 3'b110;
        rom_memory[1968] = 3'b110;
        rom_memory[1969] = 3'b110;
        rom_memory[1970] = 3'b110;
        rom_memory[1971] = 3'b110;
        rom_memory[1972] = 3'b110;
        rom_memory[1973] = 3'b110;
        rom_memory[1974] = 3'b110;
        rom_memory[1975] = 3'b110;
        rom_memory[1976] = 3'b110;
        rom_memory[1977] = 3'b110;
        rom_memory[1978] = 3'b110;
        rom_memory[1979] = 3'b110;
        rom_memory[1980] = 3'b110;
        rom_memory[1981] = 3'b110;
        rom_memory[1982] = 3'b110;
        rom_memory[1983] = 3'b110;
        rom_memory[1984] = 3'b110;
        rom_memory[1985] = 3'b110;
        rom_memory[1986] = 3'b110;
        rom_memory[1987] = 3'b110;
        rom_memory[1988] = 3'b110;
        rom_memory[1989] = 3'b110;
        rom_memory[1990] = 3'b110;
        rom_memory[1991] = 3'b110;
        rom_memory[1992] = 3'b110;
        rom_memory[1993] = 3'b110;
        rom_memory[1994] = 3'b110;
        rom_memory[1995] = 3'b110;
        rom_memory[1996] = 3'b110;
        rom_memory[1997] = 3'b110;
        rom_memory[1998] = 3'b110;
        rom_memory[1999] = 3'b110;
        rom_memory[2000] = 3'b110;
        rom_memory[2001] = 3'b110;
        rom_memory[2002] = 3'b110;
        rom_memory[2003] = 3'b110;
        rom_memory[2004] = 3'b110;
        rom_memory[2005] = 3'b110;
        rom_memory[2006] = 3'b110;
        rom_memory[2007] = 3'b110;
        rom_memory[2008] = 3'b110;
        rom_memory[2009] = 3'b110;
        rom_memory[2010] = 3'b110;
        rom_memory[2011] = 3'b110;
        rom_memory[2012] = 3'b110;
        rom_memory[2013] = 3'b110;
        rom_memory[2014] = 3'b110;
        rom_memory[2015] = 3'b110;
        rom_memory[2016] = 3'b110;
        rom_memory[2017] = 3'b110;
        rom_memory[2018] = 3'b110;
        rom_memory[2019] = 3'b110;
        rom_memory[2020] = 3'b110;
        rom_memory[2021] = 3'b110;
        rom_memory[2022] = 3'b110;
        rom_memory[2023] = 3'b110;
        rom_memory[2024] = 3'b110;
        rom_memory[2025] = 3'b110;
        rom_memory[2026] = 3'b110;
        rom_memory[2027] = 3'b110;
        rom_memory[2028] = 3'b110;
        rom_memory[2029] = 3'b110;
        rom_memory[2030] = 3'b110;
        rom_memory[2031] = 3'b110;
        rom_memory[2032] = 3'b110;
        rom_memory[2033] = 3'b110;
        rom_memory[2034] = 3'b110;
        rom_memory[2035] = 3'b110;
        rom_memory[2036] = 3'b110;
        rom_memory[2037] = 3'b110;
        rom_memory[2038] = 3'b110;
        rom_memory[2039] = 3'b110;
        rom_memory[2040] = 3'b110;
        rom_memory[2041] = 3'b110;
        rom_memory[2042] = 3'b110;
        rom_memory[2043] = 3'b110;
        rom_memory[2044] = 3'b110;
        rom_memory[2045] = 3'b110;
        rom_memory[2046] = 3'b110;
        rom_memory[2047] = 3'b110;
        rom_memory[2048] = 3'b110;
        rom_memory[2049] = 3'b110;
        rom_memory[2050] = 3'b110;
        rom_memory[2051] = 3'b110;
        rom_memory[2052] = 3'b110;
        rom_memory[2053] = 3'b110;
        rom_memory[2054] = 3'b110;
        rom_memory[2055] = 3'b110;
        rom_memory[2056] = 3'b110;
        rom_memory[2057] = 3'b110;
        rom_memory[2058] = 3'b110;
        rom_memory[2059] = 3'b110;
        rom_memory[2060] = 3'b110;
        rom_memory[2061] = 3'b110;
        rom_memory[2062] = 3'b110;
        rom_memory[2063] = 3'b110;
        rom_memory[2064] = 3'b110;
        rom_memory[2065] = 3'b110;
        rom_memory[2066] = 3'b110;
        rom_memory[2067] = 3'b110;
        rom_memory[2068] = 3'b110;
        rom_memory[2069] = 3'b110;
        rom_memory[2070] = 3'b110;
        rom_memory[2071] = 3'b110;
        rom_memory[2072] = 3'b110;
        rom_memory[2073] = 3'b110;
        rom_memory[2074] = 3'b110;
        rom_memory[2075] = 3'b110;
        rom_memory[2076] = 3'b110;
        rom_memory[2077] = 3'b110;
        rom_memory[2078] = 3'b110;
        rom_memory[2079] = 3'b110;
        rom_memory[2080] = 3'b110;
        rom_memory[2081] = 3'b100;
        rom_memory[2082] = 3'b100;
        rom_memory[2083] = 3'b100;
        rom_memory[2084] = 3'b100;
        rom_memory[2085] = 3'b100;
        rom_memory[2086] = 3'b100;
        rom_memory[2087] = 3'b100;
        rom_memory[2088] = 3'b100;
        rom_memory[2089] = 3'b100;
        rom_memory[2090] = 3'b100;
        rom_memory[2091] = 3'b100;
        rom_memory[2092] = 3'b100;
        rom_memory[2093] = 3'b100;
        rom_memory[2094] = 3'b100;
        rom_memory[2095] = 3'b100;
        rom_memory[2096] = 3'b100;
        rom_memory[2097] = 3'b100;
        rom_memory[2098] = 3'b100;
        rom_memory[2099] = 3'b100;
        rom_memory[2100] = 3'b100;
        rom_memory[2101] = 3'b100;
        rom_memory[2102] = 3'b100;
        rom_memory[2103] = 3'b100;
        rom_memory[2104] = 3'b100;
        rom_memory[2105] = 3'b100;
        rom_memory[2106] = 3'b100;
        rom_memory[2107] = 3'b100;
        rom_memory[2108] = 3'b100;
        rom_memory[2109] = 3'b100;
        rom_memory[2110] = 3'b100;
        rom_memory[2111] = 3'b100;
        rom_memory[2112] = 3'b100;
        rom_memory[2113] = 3'b100;
        rom_memory[2114] = 3'b100;
        rom_memory[2115] = 3'b100;
        rom_memory[2116] = 3'b100;
        rom_memory[2117] = 3'b100;
        rom_memory[2118] = 3'b100;
        rom_memory[2119] = 3'b100;
        rom_memory[2120] = 3'b100;
        rom_memory[2121] = 3'b100;
        rom_memory[2122] = 3'b100;
        rom_memory[2123] = 3'b100;
        rom_memory[2124] = 3'b100;
        rom_memory[2125] = 3'b100;
        rom_memory[2126] = 3'b100;
        rom_memory[2127] = 3'b100;
        rom_memory[2128] = 3'b100;
        rom_memory[2129] = 3'b100;
        rom_memory[2130] = 3'b100;
        rom_memory[2131] = 3'b100;
        rom_memory[2132] = 3'b100;
        rom_memory[2133] = 3'b100;
        rom_memory[2134] = 3'b100;
        rom_memory[2135] = 3'b100;
        rom_memory[2136] = 3'b100;
        rom_memory[2137] = 3'b100;
        rom_memory[2138] = 3'b100;
        rom_memory[2139] = 3'b100;
        rom_memory[2140] = 3'b100;
        rom_memory[2141] = 3'b100;
        rom_memory[2142] = 3'b100;
        rom_memory[2143] = 3'b100;
        rom_memory[2144] = 3'b100;
        rom_memory[2145] = 3'b100;
        rom_memory[2146] = 3'b100;
        rom_memory[2147] = 3'b100;
        rom_memory[2148] = 3'b100;
        rom_memory[2149] = 3'b100;
        rom_memory[2150] = 3'b100;
        rom_memory[2151] = 3'b100;
        rom_memory[2152] = 3'b100;
        rom_memory[2153] = 3'b100;
        rom_memory[2154] = 3'b100;
        rom_memory[2155] = 3'b100;
        rom_memory[2156] = 3'b100;
        rom_memory[2157] = 3'b100;
        rom_memory[2158] = 3'b100;
        rom_memory[2159] = 3'b100;
        rom_memory[2160] = 3'b110;
        rom_memory[2161] = 3'b110;
        rom_memory[2162] = 3'b110;
        rom_memory[2163] = 3'b110;
        rom_memory[2164] = 3'b110;
        rom_memory[2165] = 3'b110;
        rom_memory[2166] = 3'b110;
        rom_memory[2167] = 3'b110;
        rom_memory[2168] = 3'b110;
        rom_memory[2169] = 3'b110;
        rom_memory[2170] = 3'b110;
        rom_memory[2171] = 3'b110;
        rom_memory[2172] = 3'b110;
        rom_memory[2173] = 3'b110;
        rom_memory[2174] = 3'b110;
        rom_memory[2175] = 3'b110;
        rom_memory[2176] = 3'b110;
        rom_memory[2177] = 3'b110;
        rom_memory[2178] = 3'b110;
        rom_memory[2179] = 3'b110;
        rom_memory[2180] = 3'b110;
        rom_memory[2181] = 3'b110;
        rom_memory[2182] = 3'b110;
        rom_memory[2183] = 3'b110;
        rom_memory[2184] = 3'b110;
        rom_memory[2185] = 3'b110;
        rom_memory[2186] = 3'b110;
        rom_memory[2187] = 3'b110;
        rom_memory[2188] = 3'b110;
        rom_memory[2189] = 3'b110;
        rom_memory[2190] = 3'b110;
        rom_memory[2191] = 3'b110;
        rom_memory[2192] = 3'b110;
        rom_memory[2193] = 3'b110;
        rom_memory[2194] = 3'b110;
        rom_memory[2195] = 3'b110;
        rom_memory[2196] = 3'b110;
        rom_memory[2197] = 3'b110;
        rom_memory[2198] = 3'b110;
        rom_memory[2199] = 3'b110;
        rom_memory[2200] = 3'b110;
        rom_memory[2201] = 3'b110;
        rom_memory[2202] = 3'b110;
        rom_memory[2203] = 3'b110;
        rom_memory[2204] = 3'b110;
        rom_memory[2205] = 3'b110;
        rom_memory[2206] = 3'b110;
        rom_memory[2207] = 3'b110;
        rom_memory[2208] = 3'b110;
        rom_memory[2209] = 3'b110;
        rom_memory[2210] = 3'b110;
        rom_memory[2211] = 3'b110;
        rom_memory[2212] = 3'b110;
        rom_memory[2213] = 3'b110;
        rom_memory[2214] = 3'b110;
        rom_memory[2215] = 3'b110;
        rom_memory[2216] = 3'b110;
        rom_memory[2217] = 3'b110;
        rom_memory[2218] = 3'b110;
        rom_memory[2219] = 3'b110;
        rom_memory[2220] = 3'b110;
        rom_memory[2221] = 3'b110;
        rom_memory[2222] = 3'b110;
        rom_memory[2223] = 3'b110;
        rom_memory[2224] = 3'b110;
        rom_memory[2225] = 3'b110;
        rom_memory[2226] = 3'b110;
        rom_memory[2227] = 3'b110;
        rom_memory[2228] = 3'b110;
        rom_memory[2229] = 3'b110;
        rom_memory[2230] = 3'b110;
        rom_memory[2231] = 3'b110;
        rom_memory[2232] = 3'b110;
        rom_memory[2233] = 3'b110;
        rom_memory[2234] = 3'b110;
        rom_memory[2235] = 3'b110;
        rom_memory[2236] = 3'b110;
        rom_memory[2237] = 3'b110;
        rom_memory[2238] = 3'b110;
        rom_memory[2239] = 3'b110;
        rom_memory[2240] = 3'b110;
        rom_memory[2241] = 3'b110;
        rom_memory[2242] = 3'b110;
        rom_memory[2243] = 3'b110;
        rom_memory[2244] = 3'b110;
        rom_memory[2245] = 3'b110;
        rom_memory[2246] = 3'b110;
        rom_memory[2247] = 3'b110;
        rom_memory[2248] = 3'b110;
        rom_memory[2249] = 3'b110;
        rom_memory[2250] = 3'b110;
        rom_memory[2251] = 3'b110;
        rom_memory[2252] = 3'b110;
        rom_memory[2253] = 3'b110;
        rom_memory[2254] = 3'b110;
        rom_memory[2255] = 3'b110;
        rom_memory[2256] = 3'b110;
        rom_memory[2257] = 3'b110;
        rom_memory[2258] = 3'b110;
        rom_memory[2259] = 3'b110;
        rom_memory[2260] = 3'b110;
        rom_memory[2261] = 3'b110;
        rom_memory[2262] = 3'b110;
        rom_memory[2263] = 3'b110;
        rom_memory[2264] = 3'b110;
        rom_memory[2265] = 3'b110;
        rom_memory[2266] = 3'b110;
        rom_memory[2267] = 3'b110;
        rom_memory[2268] = 3'b110;
        rom_memory[2269] = 3'b110;
        rom_memory[2270] = 3'b110;
        rom_memory[2271] = 3'b110;
        rom_memory[2272] = 3'b110;
        rom_memory[2273] = 3'b110;
        rom_memory[2274] = 3'b110;
        rom_memory[2275] = 3'b110;
        rom_memory[2276] = 3'b110;
        rom_memory[2277] = 3'b110;
        rom_memory[2278] = 3'b110;
        rom_memory[2279] = 3'b110;
        rom_memory[2280] = 3'b110;
        rom_memory[2281] = 3'b110;
        rom_memory[2282] = 3'b110;
        rom_memory[2283] = 3'b110;
        rom_memory[2284] = 3'b110;
        rom_memory[2285] = 3'b110;
        rom_memory[2286] = 3'b110;
        rom_memory[2287] = 3'b110;
        rom_memory[2288] = 3'b110;
        rom_memory[2289] = 3'b110;
        rom_memory[2290] = 3'b110;
        rom_memory[2291] = 3'b110;
        rom_memory[2292] = 3'b110;
        rom_memory[2293] = 3'b110;
        rom_memory[2294] = 3'b110;
        rom_memory[2295] = 3'b110;
        rom_memory[2296] = 3'b110;
        rom_memory[2297] = 3'b110;
        rom_memory[2298] = 3'b110;
        rom_memory[2299] = 3'b110;
        rom_memory[2300] = 3'b110;
        rom_memory[2301] = 3'b110;
        rom_memory[2302] = 3'b110;
        rom_memory[2303] = 3'b110;
        rom_memory[2304] = 3'b110;
        rom_memory[2305] = 3'b110;
        rom_memory[2306] = 3'b110;
        rom_memory[2307] = 3'b110;
        rom_memory[2308] = 3'b110;
        rom_memory[2309] = 3'b110;
        rom_memory[2310] = 3'b110;
        rom_memory[2311] = 3'b110;
        rom_memory[2312] = 3'b110;
        rom_memory[2313] = 3'b110;
        rom_memory[2314] = 3'b110;
        rom_memory[2315] = 3'b110;
        rom_memory[2316] = 3'b110;
        rom_memory[2317] = 3'b110;
        rom_memory[2318] = 3'b110;
        rom_memory[2319] = 3'b110;
        rom_memory[2320] = 3'b110;
        rom_memory[2321] = 3'b110;
        rom_memory[2322] = 3'b100;
        rom_memory[2323] = 3'b100;
        rom_memory[2324] = 3'b100;
        rom_memory[2325] = 3'b100;
        rom_memory[2326] = 3'b100;
        rom_memory[2327] = 3'b100;
        rom_memory[2328] = 3'b100;
        rom_memory[2329] = 3'b100;
        rom_memory[2330] = 3'b100;
        rom_memory[2331] = 3'b100;
        rom_memory[2332] = 3'b100;
        rom_memory[2333] = 3'b100;
        rom_memory[2334] = 3'b100;
        rom_memory[2335] = 3'b100;
        rom_memory[2336] = 3'b100;
        rom_memory[2337] = 3'b100;
        rom_memory[2338] = 3'b100;
        rom_memory[2339] = 3'b100;
        rom_memory[2340] = 3'b100;
        rom_memory[2341] = 3'b100;
        rom_memory[2342] = 3'b100;
        rom_memory[2343] = 3'b100;
        rom_memory[2344] = 3'b100;
        rom_memory[2345] = 3'b100;
        rom_memory[2346] = 3'b100;
        rom_memory[2347] = 3'b100;
        rom_memory[2348] = 3'b100;
        rom_memory[2349] = 3'b100;
        rom_memory[2350] = 3'b100;
        rom_memory[2351] = 3'b100;
        rom_memory[2352] = 3'b100;
        rom_memory[2353] = 3'b100;
        rom_memory[2354] = 3'b100;
        rom_memory[2355] = 3'b100;
        rom_memory[2356] = 3'b100;
        rom_memory[2357] = 3'b100;
        rom_memory[2358] = 3'b100;
        rom_memory[2359] = 3'b100;
        rom_memory[2360] = 3'b100;
        rom_memory[2361] = 3'b100;
        rom_memory[2362] = 3'b100;
        rom_memory[2363] = 3'b100;
        rom_memory[2364] = 3'b100;
        rom_memory[2365] = 3'b100;
        rom_memory[2366] = 3'b100;
        rom_memory[2367] = 3'b100;
        rom_memory[2368] = 3'b100;
        rom_memory[2369] = 3'b100;
        rom_memory[2370] = 3'b100;
        rom_memory[2371] = 3'b100;
        rom_memory[2372] = 3'b100;
        rom_memory[2373] = 3'b100;
        rom_memory[2374] = 3'b100;
        rom_memory[2375] = 3'b100;
        rom_memory[2376] = 3'b100;
        rom_memory[2377] = 3'b100;
        rom_memory[2378] = 3'b100;
        rom_memory[2379] = 3'b100;
        rom_memory[2380] = 3'b100;
        rom_memory[2381] = 3'b100;
        rom_memory[2382] = 3'b100;
        rom_memory[2383] = 3'b100;
        rom_memory[2384] = 3'b100;
        rom_memory[2385] = 3'b100;
        rom_memory[2386] = 3'b100;
        rom_memory[2387] = 3'b100;
        rom_memory[2388] = 3'b100;
        rom_memory[2389] = 3'b100;
        rom_memory[2390] = 3'b100;
        rom_memory[2391] = 3'b100;
        rom_memory[2392] = 3'b100;
        rom_memory[2393] = 3'b100;
        rom_memory[2394] = 3'b100;
        rom_memory[2395] = 3'b100;
        rom_memory[2396] = 3'b100;
        rom_memory[2397] = 3'b100;
        rom_memory[2398] = 3'b100;
        rom_memory[2399] = 3'b100;
        rom_memory[2400] = 3'b110;
        rom_memory[2401] = 3'b110;
        rom_memory[2402] = 3'b110;
        rom_memory[2403] = 3'b110;
        rom_memory[2404] = 3'b110;
        rom_memory[2405] = 3'b110;
        rom_memory[2406] = 3'b110;
        rom_memory[2407] = 3'b110;
        rom_memory[2408] = 3'b110;
        rom_memory[2409] = 3'b110;
        rom_memory[2410] = 3'b110;
        rom_memory[2411] = 3'b110;
        rom_memory[2412] = 3'b110;
        rom_memory[2413] = 3'b110;
        rom_memory[2414] = 3'b110;
        rom_memory[2415] = 3'b110;
        rom_memory[2416] = 3'b110;
        rom_memory[2417] = 3'b110;
        rom_memory[2418] = 3'b110;
        rom_memory[2419] = 3'b110;
        rom_memory[2420] = 3'b110;
        rom_memory[2421] = 3'b110;
        rom_memory[2422] = 3'b110;
        rom_memory[2423] = 3'b110;
        rom_memory[2424] = 3'b110;
        rom_memory[2425] = 3'b110;
        rom_memory[2426] = 3'b110;
        rom_memory[2427] = 3'b110;
        rom_memory[2428] = 3'b110;
        rom_memory[2429] = 3'b110;
        rom_memory[2430] = 3'b110;
        rom_memory[2431] = 3'b110;
        rom_memory[2432] = 3'b110;
        rom_memory[2433] = 3'b110;
        rom_memory[2434] = 3'b110;
        rom_memory[2435] = 3'b110;
        rom_memory[2436] = 3'b110;
        rom_memory[2437] = 3'b110;
        rom_memory[2438] = 3'b110;
        rom_memory[2439] = 3'b110;
        rom_memory[2440] = 3'b110;
        rom_memory[2441] = 3'b110;
        rom_memory[2442] = 3'b110;
        rom_memory[2443] = 3'b110;
        rom_memory[2444] = 3'b110;
        rom_memory[2445] = 3'b110;
        rom_memory[2446] = 3'b110;
        rom_memory[2447] = 3'b110;
        rom_memory[2448] = 3'b110;
        rom_memory[2449] = 3'b110;
        rom_memory[2450] = 3'b110;
        rom_memory[2451] = 3'b110;
        rom_memory[2452] = 3'b110;
        rom_memory[2453] = 3'b110;
        rom_memory[2454] = 3'b110;
        rom_memory[2455] = 3'b110;
        rom_memory[2456] = 3'b110;
        rom_memory[2457] = 3'b110;
        rom_memory[2458] = 3'b110;
        rom_memory[2459] = 3'b110;
        rom_memory[2460] = 3'b110;
        rom_memory[2461] = 3'b110;
        rom_memory[2462] = 3'b110;
        rom_memory[2463] = 3'b110;
        rom_memory[2464] = 3'b110;
        rom_memory[2465] = 3'b110;
        rom_memory[2466] = 3'b110;
        rom_memory[2467] = 3'b110;
        rom_memory[2468] = 3'b110;
        rom_memory[2469] = 3'b110;
        rom_memory[2470] = 3'b110;
        rom_memory[2471] = 3'b110;
        rom_memory[2472] = 3'b110;
        rom_memory[2473] = 3'b110;
        rom_memory[2474] = 3'b110;
        rom_memory[2475] = 3'b110;
        rom_memory[2476] = 3'b110;
        rom_memory[2477] = 3'b110;
        rom_memory[2478] = 3'b110;
        rom_memory[2479] = 3'b110;
        rom_memory[2480] = 3'b110;
        rom_memory[2481] = 3'b110;
        rom_memory[2482] = 3'b110;
        rom_memory[2483] = 3'b110;
        rom_memory[2484] = 3'b110;
        rom_memory[2485] = 3'b110;
        rom_memory[2486] = 3'b110;
        rom_memory[2487] = 3'b110;
        rom_memory[2488] = 3'b110;
        rom_memory[2489] = 3'b110;
        rom_memory[2490] = 3'b110;
        rom_memory[2491] = 3'b110;
        rom_memory[2492] = 3'b110;
        rom_memory[2493] = 3'b110;
        rom_memory[2494] = 3'b110;
        rom_memory[2495] = 3'b110;
        rom_memory[2496] = 3'b110;
        rom_memory[2497] = 3'b110;
        rom_memory[2498] = 3'b110;
        rom_memory[2499] = 3'b110;
        rom_memory[2500] = 3'b110;
        rom_memory[2501] = 3'b110;
        rom_memory[2502] = 3'b110;
        rom_memory[2503] = 3'b110;
        rom_memory[2504] = 3'b110;
        rom_memory[2505] = 3'b110;
        rom_memory[2506] = 3'b110;
        rom_memory[2507] = 3'b110;
        rom_memory[2508] = 3'b110;
        rom_memory[2509] = 3'b110;
        rom_memory[2510] = 3'b110;
        rom_memory[2511] = 3'b110;
        rom_memory[2512] = 3'b110;
        rom_memory[2513] = 3'b110;
        rom_memory[2514] = 3'b110;
        rom_memory[2515] = 3'b110;
        rom_memory[2516] = 3'b110;
        rom_memory[2517] = 3'b110;
        rom_memory[2518] = 3'b110;
        rom_memory[2519] = 3'b110;
        rom_memory[2520] = 3'b110;
        rom_memory[2521] = 3'b110;
        rom_memory[2522] = 3'b110;
        rom_memory[2523] = 3'b110;
        rom_memory[2524] = 3'b110;
        rom_memory[2525] = 3'b110;
        rom_memory[2526] = 3'b110;
        rom_memory[2527] = 3'b110;
        rom_memory[2528] = 3'b110;
        rom_memory[2529] = 3'b110;
        rom_memory[2530] = 3'b110;
        rom_memory[2531] = 3'b110;
        rom_memory[2532] = 3'b110;
        rom_memory[2533] = 3'b110;
        rom_memory[2534] = 3'b110;
        rom_memory[2535] = 3'b110;
        rom_memory[2536] = 3'b110;
        rom_memory[2537] = 3'b110;
        rom_memory[2538] = 3'b110;
        rom_memory[2539] = 3'b110;
        rom_memory[2540] = 3'b110;
        rom_memory[2541] = 3'b110;
        rom_memory[2542] = 3'b110;
        rom_memory[2543] = 3'b110;
        rom_memory[2544] = 3'b110;
        rom_memory[2545] = 3'b110;
        rom_memory[2546] = 3'b110;
        rom_memory[2547] = 3'b110;
        rom_memory[2548] = 3'b110;
        rom_memory[2549] = 3'b110;
        rom_memory[2550] = 3'b110;
        rom_memory[2551] = 3'b110;
        rom_memory[2552] = 3'b110;
        rom_memory[2553] = 3'b110;
        rom_memory[2554] = 3'b110;
        rom_memory[2555] = 3'b110;
        rom_memory[2556] = 3'b110;
        rom_memory[2557] = 3'b110;
        rom_memory[2558] = 3'b110;
        rom_memory[2559] = 3'b110;
        rom_memory[2560] = 3'b110;
        rom_memory[2561] = 3'b110;
        rom_memory[2562] = 3'b100;
        rom_memory[2563] = 3'b100;
        rom_memory[2564] = 3'b100;
        rom_memory[2565] = 3'b100;
        rom_memory[2566] = 3'b100;
        rom_memory[2567] = 3'b100;
        rom_memory[2568] = 3'b100;
        rom_memory[2569] = 3'b100;
        rom_memory[2570] = 3'b100;
        rom_memory[2571] = 3'b100;
        rom_memory[2572] = 3'b100;
        rom_memory[2573] = 3'b100;
        rom_memory[2574] = 3'b100;
        rom_memory[2575] = 3'b100;
        rom_memory[2576] = 3'b100;
        rom_memory[2577] = 3'b100;
        rom_memory[2578] = 3'b100;
        rom_memory[2579] = 3'b100;
        rom_memory[2580] = 3'b100;
        rom_memory[2581] = 3'b100;
        rom_memory[2582] = 3'b100;
        rom_memory[2583] = 3'b100;
        rom_memory[2584] = 3'b100;
        rom_memory[2585] = 3'b100;
        rom_memory[2586] = 3'b100;
        rom_memory[2587] = 3'b100;
        rom_memory[2588] = 3'b100;
        rom_memory[2589] = 3'b100;
        rom_memory[2590] = 3'b100;
        rom_memory[2591] = 3'b100;
        rom_memory[2592] = 3'b100;
        rom_memory[2593] = 3'b100;
        rom_memory[2594] = 3'b100;
        rom_memory[2595] = 3'b100;
        rom_memory[2596] = 3'b100;
        rom_memory[2597] = 3'b100;
        rom_memory[2598] = 3'b100;
        rom_memory[2599] = 3'b100;
        rom_memory[2600] = 3'b100;
        rom_memory[2601] = 3'b100;
        rom_memory[2602] = 3'b100;
        rom_memory[2603] = 3'b100;
        rom_memory[2604] = 3'b100;
        rom_memory[2605] = 3'b100;
        rom_memory[2606] = 3'b100;
        rom_memory[2607] = 3'b100;
        rom_memory[2608] = 3'b100;
        rom_memory[2609] = 3'b100;
        rom_memory[2610] = 3'b100;
        rom_memory[2611] = 3'b100;
        rom_memory[2612] = 3'b100;
        rom_memory[2613] = 3'b100;
        rom_memory[2614] = 3'b100;
        rom_memory[2615] = 3'b100;
        rom_memory[2616] = 3'b100;
        rom_memory[2617] = 3'b100;
        rom_memory[2618] = 3'b100;
        rom_memory[2619] = 3'b100;
        rom_memory[2620] = 3'b100;
        rom_memory[2621] = 3'b100;
        rom_memory[2622] = 3'b100;
        rom_memory[2623] = 3'b100;
        rom_memory[2624] = 3'b100;
        rom_memory[2625] = 3'b100;
        rom_memory[2626] = 3'b100;
        rom_memory[2627] = 3'b100;
        rom_memory[2628] = 3'b100;
        rom_memory[2629] = 3'b100;
        rom_memory[2630] = 3'b100;
        rom_memory[2631] = 3'b100;
        rom_memory[2632] = 3'b100;
        rom_memory[2633] = 3'b100;
        rom_memory[2634] = 3'b100;
        rom_memory[2635] = 3'b100;
        rom_memory[2636] = 3'b100;
        rom_memory[2637] = 3'b100;
        rom_memory[2638] = 3'b100;
        rom_memory[2639] = 3'b100;
        rom_memory[2640] = 3'b110;
        rom_memory[2641] = 3'b110;
        rom_memory[2642] = 3'b110;
        rom_memory[2643] = 3'b110;
        rom_memory[2644] = 3'b110;
        rom_memory[2645] = 3'b110;
        rom_memory[2646] = 3'b110;
        rom_memory[2647] = 3'b110;
        rom_memory[2648] = 3'b110;
        rom_memory[2649] = 3'b110;
        rom_memory[2650] = 3'b110;
        rom_memory[2651] = 3'b110;
        rom_memory[2652] = 3'b110;
        rom_memory[2653] = 3'b110;
        rom_memory[2654] = 3'b110;
        rom_memory[2655] = 3'b110;
        rom_memory[2656] = 3'b110;
        rom_memory[2657] = 3'b110;
        rom_memory[2658] = 3'b110;
        rom_memory[2659] = 3'b110;
        rom_memory[2660] = 3'b110;
        rom_memory[2661] = 3'b110;
        rom_memory[2662] = 3'b110;
        rom_memory[2663] = 3'b110;
        rom_memory[2664] = 3'b110;
        rom_memory[2665] = 3'b110;
        rom_memory[2666] = 3'b110;
        rom_memory[2667] = 3'b110;
        rom_memory[2668] = 3'b110;
        rom_memory[2669] = 3'b110;
        rom_memory[2670] = 3'b110;
        rom_memory[2671] = 3'b110;
        rom_memory[2672] = 3'b110;
        rom_memory[2673] = 3'b110;
        rom_memory[2674] = 3'b110;
        rom_memory[2675] = 3'b110;
        rom_memory[2676] = 3'b110;
        rom_memory[2677] = 3'b110;
        rom_memory[2678] = 3'b110;
        rom_memory[2679] = 3'b110;
        rom_memory[2680] = 3'b110;
        rom_memory[2681] = 3'b110;
        rom_memory[2682] = 3'b110;
        rom_memory[2683] = 3'b110;
        rom_memory[2684] = 3'b110;
        rom_memory[2685] = 3'b110;
        rom_memory[2686] = 3'b110;
        rom_memory[2687] = 3'b110;
        rom_memory[2688] = 3'b110;
        rom_memory[2689] = 3'b110;
        rom_memory[2690] = 3'b110;
        rom_memory[2691] = 3'b110;
        rom_memory[2692] = 3'b110;
        rom_memory[2693] = 3'b110;
        rom_memory[2694] = 3'b110;
        rom_memory[2695] = 3'b110;
        rom_memory[2696] = 3'b110;
        rom_memory[2697] = 3'b110;
        rom_memory[2698] = 3'b110;
        rom_memory[2699] = 3'b110;
        rom_memory[2700] = 3'b110;
        rom_memory[2701] = 3'b110;
        rom_memory[2702] = 3'b110;
        rom_memory[2703] = 3'b110;
        rom_memory[2704] = 3'b110;
        rom_memory[2705] = 3'b110;
        rom_memory[2706] = 3'b110;
        rom_memory[2707] = 3'b110;
        rom_memory[2708] = 3'b110;
        rom_memory[2709] = 3'b110;
        rom_memory[2710] = 3'b110;
        rom_memory[2711] = 3'b110;
        rom_memory[2712] = 3'b110;
        rom_memory[2713] = 3'b110;
        rom_memory[2714] = 3'b110;
        rom_memory[2715] = 3'b110;
        rom_memory[2716] = 3'b110;
        rom_memory[2717] = 3'b110;
        rom_memory[2718] = 3'b110;
        rom_memory[2719] = 3'b110;
        rom_memory[2720] = 3'b110;
        rom_memory[2721] = 3'b110;
        rom_memory[2722] = 3'b110;
        rom_memory[2723] = 3'b110;
        rom_memory[2724] = 3'b110;
        rom_memory[2725] = 3'b110;
        rom_memory[2726] = 3'b110;
        rom_memory[2727] = 3'b110;
        rom_memory[2728] = 3'b110;
        rom_memory[2729] = 3'b110;
        rom_memory[2730] = 3'b110;
        rom_memory[2731] = 3'b110;
        rom_memory[2732] = 3'b110;
        rom_memory[2733] = 3'b110;
        rom_memory[2734] = 3'b110;
        rom_memory[2735] = 3'b110;
        rom_memory[2736] = 3'b110;
        rom_memory[2737] = 3'b110;
        rom_memory[2738] = 3'b110;
        rom_memory[2739] = 3'b110;
        rom_memory[2740] = 3'b110;
        rom_memory[2741] = 3'b110;
        rom_memory[2742] = 3'b110;
        rom_memory[2743] = 3'b110;
        rom_memory[2744] = 3'b110;
        rom_memory[2745] = 3'b110;
        rom_memory[2746] = 3'b110;
        rom_memory[2747] = 3'b110;
        rom_memory[2748] = 3'b110;
        rom_memory[2749] = 3'b110;
        rom_memory[2750] = 3'b110;
        rom_memory[2751] = 3'b110;
        rom_memory[2752] = 3'b110;
        rom_memory[2753] = 3'b110;
        rom_memory[2754] = 3'b110;
        rom_memory[2755] = 3'b110;
        rom_memory[2756] = 3'b110;
        rom_memory[2757] = 3'b110;
        rom_memory[2758] = 3'b110;
        rom_memory[2759] = 3'b110;
        rom_memory[2760] = 3'b110;
        rom_memory[2761] = 3'b110;
        rom_memory[2762] = 3'b110;
        rom_memory[2763] = 3'b110;
        rom_memory[2764] = 3'b110;
        rom_memory[2765] = 3'b110;
        rom_memory[2766] = 3'b110;
        rom_memory[2767] = 3'b110;
        rom_memory[2768] = 3'b110;
        rom_memory[2769] = 3'b110;
        rom_memory[2770] = 3'b110;
        rom_memory[2771] = 3'b110;
        rom_memory[2772] = 3'b110;
        rom_memory[2773] = 3'b110;
        rom_memory[2774] = 3'b110;
        rom_memory[2775] = 3'b110;
        rom_memory[2776] = 3'b110;
        rom_memory[2777] = 3'b110;
        rom_memory[2778] = 3'b110;
        rom_memory[2779] = 3'b110;
        rom_memory[2780] = 3'b110;
        rom_memory[2781] = 3'b110;
        rom_memory[2782] = 3'b110;
        rom_memory[2783] = 3'b110;
        rom_memory[2784] = 3'b110;
        rom_memory[2785] = 3'b110;
        rom_memory[2786] = 3'b110;
        rom_memory[2787] = 3'b110;
        rom_memory[2788] = 3'b110;
        rom_memory[2789] = 3'b110;
        rom_memory[2790] = 3'b110;
        rom_memory[2791] = 3'b110;
        rom_memory[2792] = 3'b110;
        rom_memory[2793] = 3'b110;
        rom_memory[2794] = 3'b110;
        rom_memory[2795] = 3'b110;
        rom_memory[2796] = 3'b110;
        rom_memory[2797] = 3'b110;
        rom_memory[2798] = 3'b110;
        rom_memory[2799] = 3'b110;
        rom_memory[2800] = 3'b110;
        rom_memory[2801] = 3'b110;
        rom_memory[2802] = 3'b100;
        rom_memory[2803] = 3'b100;
        rom_memory[2804] = 3'b100;
        rom_memory[2805] = 3'b100;
        rom_memory[2806] = 3'b100;
        rom_memory[2807] = 3'b100;
        rom_memory[2808] = 3'b100;
        rom_memory[2809] = 3'b100;
        rom_memory[2810] = 3'b100;
        rom_memory[2811] = 3'b100;
        rom_memory[2812] = 3'b100;
        rom_memory[2813] = 3'b100;
        rom_memory[2814] = 3'b100;
        rom_memory[2815] = 3'b100;
        rom_memory[2816] = 3'b100;
        rom_memory[2817] = 3'b100;
        rom_memory[2818] = 3'b100;
        rom_memory[2819] = 3'b100;
        rom_memory[2820] = 3'b100;
        rom_memory[2821] = 3'b100;
        rom_memory[2822] = 3'b100;
        rom_memory[2823] = 3'b100;
        rom_memory[2824] = 3'b100;
        rom_memory[2825] = 3'b100;
        rom_memory[2826] = 3'b100;
        rom_memory[2827] = 3'b100;
        rom_memory[2828] = 3'b100;
        rom_memory[2829] = 3'b100;
        rom_memory[2830] = 3'b100;
        rom_memory[2831] = 3'b100;
        rom_memory[2832] = 3'b100;
        rom_memory[2833] = 3'b100;
        rom_memory[2834] = 3'b100;
        rom_memory[2835] = 3'b100;
        rom_memory[2836] = 3'b100;
        rom_memory[2837] = 3'b100;
        rom_memory[2838] = 3'b100;
        rom_memory[2839] = 3'b100;
        rom_memory[2840] = 3'b100;
        rom_memory[2841] = 3'b100;
        rom_memory[2842] = 3'b100;
        rom_memory[2843] = 3'b100;
        rom_memory[2844] = 3'b100;
        rom_memory[2845] = 3'b100;
        rom_memory[2846] = 3'b100;
        rom_memory[2847] = 3'b100;
        rom_memory[2848] = 3'b100;
        rom_memory[2849] = 3'b100;
        rom_memory[2850] = 3'b100;
        rom_memory[2851] = 3'b100;
        rom_memory[2852] = 3'b100;
        rom_memory[2853] = 3'b100;
        rom_memory[2854] = 3'b100;
        rom_memory[2855] = 3'b100;
        rom_memory[2856] = 3'b100;
        rom_memory[2857] = 3'b100;
        rom_memory[2858] = 3'b100;
        rom_memory[2859] = 3'b100;
        rom_memory[2860] = 3'b100;
        rom_memory[2861] = 3'b100;
        rom_memory[2862] = 3'b100;
        rom_memory[2863] = 3'b100;
        rom_memory[2864] = 3'b100;
        rom_memory[2865] = 3'b100;
        rom_memory[2866] = 3'b100;
        rom_memory[2867] = 3'b100;
        rom_memory[2868] = 3'b100;
        rom_memory[2869] = 3'b100;
        rom_memory[2870] = 3'b100;
        rom_memory[2871] = 3'b100;
        rom_memory[2872] = 3'b100;
        rom_memory[2873] = 3'b100;
        rom_memory[2874] = 3'b100;
        rom_memory[2875] = 3'b100;
        rom_memory[2876] = 3'b100;
        rom_memory[2877] = 3'b100;
        rom_memory[2878] = 3'b100;
        rom_memory[2879] = 3'b100;
        rom_memory[2880] = 3'b110;
        rom_memory[2881] = 3'b110;
        rom_memory[2882] = 3'b110;
        rom_memory[2883] = 3'b110;
        rom_memory[2884] = 3'b110;
        rom_memory[2885] = 3'b110;
        rom_memory[2886] = 3'b110;
        rom_memory[2887] = 3'b110;
        rom_memory[2888] = 3'b110;
        rom_memory[2889] = 3'b110;
        rom_memory[2890] = 3'b110;
        rom_memory[2891] = 3'b110;
        rom_memory[2892] = 3'b110;
        rom_memory[2893] = 3'b110;
        rom_memory[2894] = 3'b110;
        rom_memory[2895] = 3'b110;
        rom_memory[2896] = 3'b110;
        rom_memory[2897] = 3'b110;
        rom_memory[2898] = 3'b110;
        rom_memory[2899] = 3'b110;
        rom_memory[2900] = 3'b110;
        rom_memory[2901] = 3'b110;
        rom_memory[2902] = 3'b110;
        rom_memory[2903] = 3'b110;
        rom_memory[2904] = 3'b110;
        rom_memory[2905] = 3'b110;
        rom_memory[2906] = 3'b110;
        rom_memory[2907] = 3'b110;
        rom_memory[2908] = 3'b110;
        rom_memory[2909] = 3'b110;
        rom_memory[2910] = 3'b110;
        rom_memory[2911] = 3'b110;
        rom_memory[2912] = 3'b110;
        rom_memory[2913] = 3'b110;
        rom_memory[2914] = 3'b110;
        rom_memory[2915] = 3'b110;
        rom_memory[2916] = 3'b110;
        rom_memory[2917] = 3'b110;
        rom_memory[2918] = 3'b110;
        rom_memory[2919] = 3'b110;
        rom_memory[2920] = 3'b110;
        rom_memory[2921] = 3'b110;
        rom_memory[2922] = 3'b110;
        rom_memory[2923] = 3'b110;
        rom_memory[2924] = 3'b110;
        rom_memory[2925] = 3'b110;
        rom_memory[2926] = 3'b110;
        rom_memory[2927] = 3'b110;
        rom_memory[2928] = 3'b110;
        rom_memory[2929] = 3'b110;
        rom_memory[2930] = 3'b110;
        rom_memory[2931] = 3'b110;
        rom_memory[2932] = 3'b110;
        rom_memory[2933] = 3'b110;
        rom_memory[2934] = 3'b110;
        rom_memory[2935] = 3'b110;
        rom_memory[2936] = 3'b110;
        rom_memory[2937] = 3'b110;
        rom_memory[2938] = 3'b110;
        rom_memory[2939] = 3'b110;
        rom_memory[2940] = 3'b110;
        rom_memory[2941] = 3'b110;
        rom_memory[2942] = 3'b110;
        rom_memory[2943] = 3'b110;
        rom_memory[2944] = 3'b110;
        rom_memory[2945] = 3'b110;
        rom_memory[2946] = 3'b110;
        rom_memory[2947] = 3'b110;
        rom_memory[2948] = 3'b110;
        rom_memory[2949] = 3'b110;
        rom_memory[2950] = 3'b110;
        rom_memory[2951] = 3'b110;
        rom_memory[2952] = 3'b110;
        rom_memory[2953] = 3'b110;
        rom_memory[2954] = 3'b110;
        rom_memory[2955] = 3'b110;
        rom_memory[2956] = 3'b110;
        rom_memory[2957] = 3'b110;
        rom_memory[2958] = 3'b110;
        rom_memory[2959] = 3'b110;
        rom_memory[2960] = 3'b110;
        rom_memory[2961] = 3'b110;
        rom_memory[2962] = 3'b110;
        rom_memory[2963] = 3'b110;
        rom_memory[2964] = 3'b110;
        rom_memory[2965] = 3'b110;
        rom_memory[2966] = 3'b110;
        rom_memory[2967] = 3'b110;
        rom_memory[2968] = 3'b110;
        rom_memory[2969] = 3'b110;
        rom_memory[2970] = 3'b110;
        rom_memory[2971] = 3'b110;
        rom_memory[2972] = 3'b110;
        rom_memory[2973] = 3'b110;
        rom_memory[2974] = 3'b110;
        rom_memory[2975] = 3'b110;
        rom_memory[2976] = 3'b110;
        rom_memory[2977] = 3'b110;
        rom_memory[2978] = 3'b110;
        rom_memory[2979] = 3'b110;
        rom_memory[2980] = 3'b110;
        rom_memory[2981] = 3'b110;
        rom_memory[2982] = 3'b110;
        rom_memory[2983] = 3'b110;
        rom_memory[2984] = 3'b110;
        rom_memory[2985] = 3'b110;
        rom_memory[2986] = 3'b110;
        rom_memory[2987] = 3'b110;
        rom_memory[2988] = 3'b110;
        rom_memory[2989] = 3'b110;
        rom_memory[2990] = 3'b110;
        rom_memory[2991] = 3'b110;
        rom_memory[2992] = 3'b110;
        rom_memory[2993] = 3'b110;
        rom_memory[2994] = 3'b110;
        rom_memory[2995] = 3'b110;
        rom_memory[2996] = 3'b110;
        rom_memory[2997] = 3'b110;
        rom_memory[2998] = 3'b110;
        rom_memory[2999] = 3'b110;
        rom_memory[3000] = 3'b110;
        rom_memory[3001] = 3'b110;
        rom_memory[3002] = 3'b110;
        rom_memory[3003] = 3'b110;
        rom_memory[3004] = 3'b110;
        rom_memory[3005] = 3'b110;
        rom_memory[3006] = 3'b110;
        rom_memory[3007] = 3'b110;
        rom_memory[3008] = 3'b110;
        rom_memory[3009] = 3'b110;
        rom_memory[3010] = 3'b110;
        rom_memory[3011] = 3'b110;
        rom_memory[3012] = 3'b110;
        rom_memory[3013] = 3'b110;
        rom_memory[3014] = 3'b110;
        rom_memory[3015] = 3'b110;
        rom_memory[3016] = 3'b110;
        rom_memory[3017] = 3'b110;
        rom_memory[3018] = 3'b110;
        rom_memory[3019] = 3'b110;
        rom_memory[3020] = 3'b110;
        rom_memory[3021] = 3'b110;
        rom_memory[3022] = 3'b110;
        rom_memory[3023] = 3'b110;
        rom_memory[3024] = 3'b110;
        rom_memory[3025] = 3'b110;
        rom_memory[3026] = 3'b110;
        rom_memory[3027] = 3'b110;
        rom_memory[3028] = 3'b110;
        rom_memory[3029] = 3'b110;
        rom_memory[3030] = 3'b110;
        rom_memory[3031] = 3'b110;
        rom_memory[3032] = 3'b110;
        rom_memory[3033] = 3'b110;
        rom_memory[3034] = 3'b110;
        rom_memory[3035] = 3'b110;
        rom_memory[3036] = 3'b110;
        rom_memory[3037] = 3'b110;
        rom_memory[3038] = 3'b110;
        rom_memory[3039] = 3'b110;
        rom_memory[3040] = 3'b110;
        rom_memory[3041] = 3'b110;
        rom_memory[3042] = 3'b100;
        rom_memory[3043] = 3'b100;
        rom_memory[3044] = 3'b100;
        rom_memory[3045] = 3'b100;
        rom_memory[3046] = 3'b100;
        rom_memory[3047] = 3'b100;
        rom_memory[3048] = 3'b100;
        rom_memory[3049] = 3'b100;
        rom_memory[3050] = 3'b100;
        rom_memory[3051] = 3'b100;
        rom_memory[3052] = 3'b100;
        rom_memory[3053] = 3'b100;
        rom_memory[3054] = 3'b100;
        rom_memory[3055] = 3'b100;
        rom_memory[3056] = 3'b100;
        rom_memory[3057] = 3'b100;
        rom_memory[3058] = 3'b100;
        rom_memory[3059] = 3'b100;
        rom_memory[3060] = 3'b100;
        rom_memory[3061] = 3'b100;
        rom_memory[3062] = 3'b100;
        rom_memory[3063] = 3'b100;
        rom_memory[3064] = 3'b100;
        rom_memory[3065] = 3'b100;
        rom_memory[3066] = 3'b100;
        rom_memory[3067] = 3'b100;
        rom_memory[3068] = 3'b100;
        rom_memory[3069] = 3'b100;
        rom_memory[3070] = 3'b100;
        rom_memory[3071] = 3'b100;
        rom_memory[3072] = 3'b100;
        rom_memory[3073] = 3'b100;
        rom_memory[3074] = 3'b100;
        rom_memory[3075] = 3'b100;
        rom_memory[3076] = 3'b100;
        rom_memory[3077] = 3'b100;
        rom_memory[3078] = 3'b100;
        rom_memory[3079] = 3'b100;
        rom_memory[3080] = 3'b100;
        rom_memory[3081] = 3'b100;
        rom_memory[3082] = 3'b100;
        rom_memory[3083] = 3'b100;
        rom_memory[3084] = 3'b100;
        rom_memory[3085] = 3'b100;
        rom_memory[3086] = 3'b100;
        rom_memory[3087] = 3'b100;
        rom_memory[3088] = 3'b100;
        rom_memory[3089] = 3'b100;
        rom_memory[3090] = 3'b100;
        rom_memory[3091] = 3'b100;
        rom_memory[3092] = 3'b100;
        rom_memory[3093] = 3'b100;
        rom_memory[3094] = 3'b100;
        rom_memory[3095] = 3'b100;
        rom_memory[3096] = 3'b100;
        rom_memory[3097] = 3'b100;
        rom_memory[3098] = 3'b100;
        rom_memory[3099] = 3'b100;
        rom_memory[3100] = 3'b100;
        rom_memory[3101] = 3'b100;
        rom_memory[3102] = 3'b100;
        rom_memory[3103] = 3'b100;
        rom_memory[3104] = 3'b100;
        rom_memory[3105] = 3'b100;
        rom_memory[3106] = 3'b100;
        rom_memory[3107] = 3'b100;
        rom_memory[3108] = 3'b100;
        rom_memory[3109] = 3'b100;
        rom_memory[3110] = 3'b100;
        rom_memory[3111] = 3'b110;
        rom_memory[3112] = 3'b100;
        rom_memory[3113] = 3'b100;
        rom_memory[3114] = 3'b110;
        rom_memory[3115] = 3'b100;
        rom_memory[3116] = 3'b100;
        rom_memory[3117] = 3'b100;
        rom_memory[3118] = 3'b100;
        rom_memory[3119] = 3'b100;
        rom_memory[3120] = 3'b110;
        rom_memory[3121] = 3'b110;
        rom_memory[3122] = 3'b110;
        rom_memory[3123] = 3'b110;
        rom_memory[3124] = 3'b110;
        rom_memory[3125] = 3'b110;
        rom_memory[3126] = 3'b110;
        rom_memory[3127] = 3'b110;
        rom_memory[3128] = 3'b110;
        rom_memory[3129] = 3'b110;
        rom_memory[3130] = 3'b110;
        rom_memory[3131] = 3'b110;
        rom_memory[3132] = 3'b110;
        rom_memory[3133] = 3'b110;
        rom_memory[3134] = 3'b110;
        rom_memory[3135] = 3'b110;
        rom_memory[3136] = 3'b110;
        rom_memory[3137] = 3'b110;
        rom_memory[3138] = 3'b110;
        rom_memory[3139] = 3'b110;
        rom_memory[3140] = 3'b110;
        rom_memory[3141] = 3'b110;
        rom_memory[3142] = 3'b110;
        rom_memory[3143] = 3'b110;
        rom_memory[3144] = 3'b110;
        rom_memory[3145] = 3'b110;
        rom_memory[3146] = 3'b110;
        rom_memory[3147] = 3'b110;
        rom_memory[3148] = 3'b110;
        rom_memory[3149] = 3'b110;
        rom_memory[3150] = 3'b110;
        rom_memory[3151] = 3'b110;
        rom_memory[3152] = 3'b110;
        rom_memory[3153] = 3'b110;
        rom_memory[3154] = 3'b110;
        rom_memory[3155] = 3'b110;
        rom_memory[3156] = 3'b110;
        rom_memory[3157] = 3'b110;
        rom_memory[3158] = 3'b110;
        rom_memory[3159] = 3'b110;
        rom_memory[3160] = 3'b110;
        rom_memory[3161] = 3'b110;
        rom_memory[3162] = 3'b110;
        rom_memory[3163] = 3'b110;
        rom_memory[3164] = 3'b110;
        rom_memory[3165] = 3'b110;
        rom_memory[3166] = 3'b110;
        rom_memory[3167] = 3'b110;
        rom_memory[3168] = 3'b110;
        rom_memory[3169] = 3'b110;
        rom_memory[3170] = 3'b110;
        rom_memory[3171] = 3'b110;
        rom_memory[3172] = 3'b110;
        rom_memory[3173] = 3'b110;
        rom_memory[3174] = 3'b110;
        rom_memory[3175] = 3'b110;
        rom_memory[3176] = 3'b110;
        rom_memory[3177] = 3'b110;
        rom_memory[3178] = 3'b110;
        rom_memory[3179] = 3'b110;
        rom_memory[3180] = 3'b110;
        rom_memory[3181] = 3'b110;
        rom_memory[3182] = 3'b110;
        rom_memory[3183] = 3'b110;
        rom_memory[3184] = 3'b110;
        rom_memory[3185] = 3'b110;
        rom_memory[3186] = 3'b110;
        rom_memory[3187] = 3'b110;
        rom_memory[3188] = 3'b110;
        rom_memory[3189] = 3'b110;
        rom_memory[3190] = 3'b110;
        rom_memory[3191] = 3'b110;
        rom_memory[3192] = 3'b110;
        rom_memory[3193] = 3'b110;
        rom_memory[3194] = 3'b110;
        rom_memory[3195] = 3'b110;
        rom_memory[3196] = 3'b110;
        rom_memory[3197] = 3'b110;
        rom_memory[3198] = 3'b110;
        rom_memory[3199] = 3'b110;
        rom_memory[3200] = 3'b110;
        rom_memory[3201] = 3'b110;
        rom_memory[3202] = 3'b110;
        rom_memory[3203] = 3'b110;
        rom_memory[3204] = 3'b110;
        rom_memory[3205] = 3'b110;
        rom_memory[3206] = 3'b110;
        rom_memory[3207] = 3'b110;
        rom_memory[3208] = 3'b110;
        rom_memory[3209] = 3'b110;
        rom_memory[3210] = 3'b110;
        rom_memory[3211] = 3'b110;
        rom_memory[3212] = 3'b110;
        rom_memory[3213] = 3'b110;
        rom_memory[3214] = 3'b110;
        rom_memory[3215] = 3'b110;
        rom_memory[3216] = 3'b110;
        rom_memory[3217] = 3'b110;
        rom_memory[3218] = 3'b110;
        rom_memory[3219] = 3'b110;
        rom_memory[3220] = 3'b110;
        rom_memory[3221] = 3'b110;
        rom_memory[3222] = 3'b110;
        rom_memory[3223] = 3'b110;
        rom_memory[3224] = 3'b110;
        rom_memory[3225] = 3'b110;
        rom_memory[3226] = 3'b110;
        rom_memory[3227] = 3'b110;
        rom_memory[3228] = 3'b110;
        rom_memory[3229] = 3'b110;
        rom_memory[3230] = 3'b110;
        rom_memory[3231] = 3'b110;
        rom_memory[3232] = 3'b110;
        rom_memory[3233] = 3'b110;
        rom_memory[3234] = 3'b110;
        rom_memory[3235] = 3'b110;
        rom_memory[3236] = 3'b110;
        rom_memory[3237] = 3'b110;
        rom_memory[3238] = 3'b110;
        rom_memory[3239] = 3'b110;
        rom_memory[3240] = 3'b110;
        rom_memory[3241] = 3'b110;
        rom_memory[3242] = 3'b110;
        rom_memory[3243] = 3'b110;
        rom_memory[3244] = 3'b110;
        rom_memory[3245] = 3'b110;
        rom_memory[3246] = 3'b110;
        rom_memory[3247] = 3'b110;
        rom_memory[3248] = 3'b110;
        rom_memory[3249] = 3'b110;
        rom_memory[3250] = 3'b110;
        rom_memory[3251] = 3'b110;
        rom_memory[3252] = 3'b110;
        rom_memory[3253] = 3'b110;
        rom_memory[3254] = 3'b110;
        rom_memory[3255] = 3'b110;
        rom_memory[3256] = 3'b110;
        rom_memory[3257] = 3'b110;
        rom_memory[3258] = 3'b110;
        rom_memory[3259] = 3'b110;
        rom_memory[3260] = 3'b110;
        rom_memory[3261] = 3'b110;
        rom_memory[3262] = 3'b110;
        rom_memory[3263] = 3'b110;
        rom_memory[3264] = 3'b110;
        rom_memory[3265] = 3'b110;
        rom_memory[3266] = 3'b110;
        rom_memory[3267] = 3'b110;
        rom_memory[3268] = 3'b110;
        rom_memory[3269] = 3'b110;
        rom_memory[3270] = 3'b110;
        rom_memory[3271] = 3'b110;
        rom_memory[3272] = 3'b110;
        rom_memory[3273] = 3'b110;
        rom_memory[3274] = 3'b110;
        rom_memory[3275] = 3'b110;
        rom_memory[3276] = 3'b110;
        rom_memory[3277] = 3'b110;
        rom_memory[3278] = 3'b110;
        rom_memory[3279] = 3'b110;
        rom_memory[3280] = 3'b110;
        rom_memory[3281] = 3'b110;
        rom_memory[3282] = 3'b110;
        rom_memory[3283] = 3'b110;
        rom_memory[3284] = 3'b110;
        rom_memory[3285] = 3'b110;
        rom_memory[3286] = 3'b110;
        rom_memory[3287] = 3'b100;
        rom_memory[3288] = 3'b100;
        rom_memory[3289] = 3'b100;
        rom_memory[3290] = 3'b100;
        rom_memory[3291] = 3'b100;
        rom_memory[3292] = 3'b100;
        rom_memory[3293] = 3'b100;
        rom_memory[3294] = 3'b100;
        rom_memory[3295] = 3'b100;
        rom_memory[3296] = 3'b100;
        rom_memory[3297] = 3'b100;
        rom_memory[3298] = 3'b100;
        rom_memory[3299] = 3'b100;
        rom_memory[3300] = 3'b100;
        rom_memory[3301] = 3'b100;
        rom_memory[3302] = 3'b100;
        rom_memory[3303] = 3'b100;
        rom_memory[3304] = 3'b100;
        rom_memory[3305] = 3'b100;
        rom_memory[3306] = 3'b100;
        rom_memory[3307] = 3'b100;
        rom_memory[3308] = 3'b100;
        rom_memory[3309] = 3'b100;
        rom_memory[3310] = 3'b100;
        rom_memory[3311] = 3'b100;
        rom_memory[3312] = 3'b100;
        rom_memory[3313] = 3'b100;
        rom_memory[3314] = 3'b100;
        rom_memory[3315] = 3'b100;
        rom_memory[3316] = 3'b100;
        rom_memory[3317] = 3'b100;
        rom_memory[3318] = 3'b100;
        rom_memory[3319] = 3'b100;
        rom_memory[3320] = 3'b100;
        rom_memory[3321] = 3'b100;
        rom_memory[3322] = 3'b100;
        rom_memory[3323] = 3'b100;
        rom_memory[3324] = 3'b100;
        rom_memory[3325] = 3'b100;
        rom_memory[3326] = 3'b100;
        rom_memory[3327] = 3'b100;
        rom_memory[3328] = 3'b100;
        rom_memory[3329] = 3'b100;
        rom_memory[3330] = 3'b100;
        rom_memory[3331] = 3'b100;
        rom_memory[3332] = 3'b100;
        rom_memory[3333] = 3'b100;
        rom_memory[3334] = 3'b100;
        rom_memory[3335] = 3'b100;
        rom_memory[3336] = 3'b100;
        rom_memory[3337] = 3'b100;
        rom_memory[3338] = 3'b100;
        rom_memory[3339] = 3'b100;
        rom_memory[3340] = 3'b100;
        rom_memory[3341] = 3'b100;
        rom_memory[3342] = 3'b100;
        rom_memory[3343] = 3'b100;
        rom_memory[3344] = 3'b100;
        rom_memory[3345] = 3'b100;
        rom_memory[3346] = 3'b110;
        rom_memory[3347] = 3'b100;
        rom_memory[3348] = 3'b100;
        rom_memory[3349] = 3'b100;
        rom_memory[3350] = 3'b100;
        rom_memory[3351] = 3'b100;
        rom_memory[3352] = 3'b100;
        rom_memory[3353] = 3'b100;
        rom_memory[3354] = 3'b100;
        rom_memory[3355] = 3'b110;
        rom_memory[3356] = 3'b100;
        rom_memory[3357] = 3'b100;
        rom_memory[3358] = 3'b110;
        rom_memory[3359] = 3'b110;
        rom_memory[3360] = 3'b110;
        rom_memory[3361] = 3'b110;
        rom_memory[3362] = 3'b110;
        rom_memory[3363] = 3'b110;
        rom_memory[3364] = 3'b110;
        rom_memory[3365] = 3'b110;
        rom_memory[3366] = 3'b110;
        rom_memory[3367] = 3'b110;
        rom_memory[3368] = 3'b110;
        rom_memory[3369] = 3'b110;
        rom_memory[3370] = 3'b110;
        rom_memory[3371] = 3'b110;
        rom_memory[3372] = 3'b110;
        rom_memory[3373] = 3'b110;
        rom_memory[3374] = 3'b110;
        rom_memory[3375] = 3'b110;
        rom_memory[3376] = 3'b110;
        rom_memory[3377] = 3'b110;
        rom_memory[3378] = 3'b110;
        rom_memory[3379] = 3'b110;
        rom_memory[3380] = 3'b110;
        rom_memory[3381] = 3'b110;
        rom_memory[3382] = 3'b110;
        rom_memory[3383] = 3'b110;
        rom_memory[3384] = 3'b110;
        rom_memory[3385] = 3'b110;
        rom_memory[3386] = 3'b110;
        rom_memory[3387] = 3'b110;
        rom_memory[3388] = 3'b110;
        rom_memory[3389] = 3'b110;
        rom_memory[3390] = 3'b110;
        rom_memory[3391] = 3'b110;
        rom_memory[3392] = 3'b110;
        rom_memory[3393] = 3'b110;
        rom_memory[3394] = 3'b110;
        rom_memory[3395] = 3'b110;
        rom_memory[3396] = 3'b110;
        rom_memory[3397] = 3'b110;
        rom_memory[3398] = 3'b110;
        rom_memory[3399] = 3'b110;
        rom_memory[3400] = 3'b110;
        rom_memory[3401] = 3'b110;
        rom_memory[3402] = 3'b110;
        rom_memory[3403] = 3'b110;
        rom_memory[3404] = 3'b110;
        rom_memory[3405] = 3'b110;
        rom_memory[3406] = 3'b110;
        rom_memory[3407] = 3'b110;
        rom_memory[3408] = 3'b110;
        rom_memory[3409] = 3'b110;
        rom_memory[3410] = 3'b110;
        rom_memory[3411] = 3'b110;
        rom_memory[3412] = 3'b110;
        rom_memory[3413] = 3'b110;
        rom_memory[3414] = 3'b110;
        rom_memory[3415] = 3'b110;
        rom_memory[3416] = 3'b110;
        rom_memory[3417] = 3'b110;
        rom_memory[3418] = 3'b110;
        rom_memory[3419] = 3'b110;
        rom_memory[3420] = 3'b110;
        rom_memory[3421] = 3'b110;
        rom_memory[3422] = 3'b110;
        rom_memory[3423] = 3'b110;
        rom_memory[3424] = 3'b110;
        rom_memory[3425] = 3'b110;
        rom_memory[3426] = 3'b110;
        rom_memory[3427] = 3'b110;
        rom_memory[3428] = 3'b110;
        rom_memory[3429] = 3'b110;
        rom_memory[3430] = 3'b110;
        rom_memory[3431] = 3'b110;
        rom_memory[3432] = 3'b110;
        rom_memory[3433] = 3'b110;
        rom_memory[3434] = 3'b110;
        rom_memory[3435] = 3'b110;
        rom_memory[3436] = 3'b110;
        rom_memory[3437] = 3'b110;
        rom_memory[3438] = 3'b110;
        rom_memory[3439] = 3'b110;
        rom_memory[3440] = 3'b110;
        rom_memory[3441] = 3'b110;
        rom_memory[3442] = 3'b110;
        rom_memory[3443] = 3'b110;
        rom_memory[3444] = 3'b110;
        rom_memory[3445] = 3'b110;
        rom_memory[3446] = 3'b110;
        rom_memory[3447] = 3'b110;
        rom_memory[3448] = 3'b110;
        rom_memory[3449] = 3'b110;
        rom_memory[3450] = 3'b110;
        rom_memory[3451] = 3'b110;
        rom_memory[3452] = 3'b110;
        rom_memory[3453] = 3'b110;
        rom_memory[3454] = 3'b110;
        rom_memory[3455] = 3'b110;
        rom_memory[3456] = 3'b110;
        rom_memory[3457] = 3'b110;
        rom_memory[3458] = 3'b110;
        rom_memory[3459] = 3'b110;
        rom_memory[3460] = 3'b110;
        rom_memory[3461] = 3'b110;
        rom_memory[3462] = 3'b110;
        rom_memory[3463] = 3'b110;
        rom_memory[3464] = 3'b110;
        rom_memory[3465] = 3'b110;
        rom_memory[3466] = 3'b110;
        rom_memory[3467] = 3'b110;
        rom_memory[3468] = 3'b110;
        rom_memory[3469] = 3'b110;
        rom_memory[3470] = 3'b110;
        rom_memory[3471] = 3'b110;
        rom_memory[3472] = 3'b110;
        rom_memory[3473] = 3'b110;
        rom_memory[3474] = 3'b110;
        rom_memory[3475] = 3'b110;
        rom_memory[3476] = 3'b110;
        rom_memory[3477] = 3'b110;
        rom_memory[3478] = 3'b110;
        rom_memory[3479] = 3'b110;
        rom_memory[3480] = 3'b110;
        rom_memory[3481] = 3'b110;
        rom_memory[3482] = 3'b110;
        rom_memory[3483] = 3'b110;
        rom_memory[3484] = 3'b110;
        rom_memory[3485] = 3'b110;
        rom_memory[3486] = 3'b110;
        rom_memory[3487] = 3'b110;
        rom_memory[3488] = 3'b110;
        rom_memory[3489] = 3'b110;
        rom_memory[3490] = 3'b110;
        rom_memory[3491] = 3'b110;
        rom_memory[3492] = 3'b110;
        rom_memory[3493] = 3'b110;
        rom_memory[3494] = 3'b110;
        rom_memory[3495] = 3'b110;
        rom_memory[3496] = 3'b110;
        rom_memory[3497] = 3'b110;
        rom_memory[3498] = 3'b110;
        rom_memory[3499] = 3'b110;
        rom_memory[3500] = 3'b110;
        rom_memory[3501] = 3'b110;
        rom_memory[3502] = 3'b110;
        rom_memory[3503] = 3'b110;
        rom_memory[3504] = 3'b110;
        rom_memory[3505] = 3'b110;
        rom_memory[3506] = 3'b110;
        rom_memory[3507] = 3'b110;
        rom_memory[3508] = 3'b110;
        rom_memory[3509] = 3'b110;
        rom_memory[3510] = 3'b110;
        rom_memory[3511] = 3'b110;
        rom_memory[3512] = 3'b110;
        rom_memory[3513] = 3'b110;
        rom_memory[3514] = 3'b110;
        rom_memory[3515] = 3'b110;
        rom_memory[3516] = 3'b110;
        rom_memory[3517] = 3'b110;
        rom_memory[3518] = 3'b110;
        rom_memory[3519] = 3'b110;
        rom_memory[3520] = 3'b110;
        rom_memory[3521] = 3'b110;
        rom_memory[3522] = 3'b110;
        rom_memory[3523] = 3'b110;
        rom_memory[3524] = 3'b110;
        rom_memory[3525] = 3'b110;
        rom_memory[3526] = 3'b110;
        rom_memory[3527] = 3'b110;
        rom_memory[3528] = 3'b100;
        rom_memory[3529] = 3'b100;
        rom_memory[3530] = 3'b100;
        rom_memory[3531] = 3'b100;
        rom_memory[3532] = 3'b110;
        rom_memory[3533] = 3'b100;
        rom_memory[3534] = 3'b100;
        rom_memory[3535] = 3'b100;
        rom_memory[3536] = 3'b100;
        rom_memory[3537] = 3'b100;
        rom_memory[3538] = 3'b100;
        rom_memory[3539] = 3'b100;
        rom_memory[3540] = 3'b100;
        rom_memory[3541] = 3'b100;
        rom_memory[3542] = 3'b100;
        rom_memory[3543] = 3'b100;
        rom_memory[3544] = 3'b100;
        rom_memory[3545] = 3'b100;
        rom_memory[3546] = 3'b100;
        rom_memory[3547] = 3'b100;
        rom_memory[3548] = 3'b100;
        rom_memory[3549] = 3'b100;
        rom_memory[3550] = 3'b100;
        rom_memory[3551] = 3'b100;
        rom_memory[3552] = 3'b100;
        rom_memory[3553] = 3'b110;
        rom_memory[3554] = 3'b110;
        rom_memory[3555] = 3'b100;
        rom_memory[3556] = 3'b100;
        rom_memory[3557] = 3'b100;
        rom_memory[3558] = 3'b100;
        rom_memory[3559] = 3'b100;
        rom_memory[3560] = 3'b110;
        rom_memory[3561] = 3'b100;
        rom_memory[3562] = 3'b100;
        rom_memory[3563] = 3'b100;
        rom_memory[3564] = 3'b100;
        rom_memory[3565] = 3'b100;
        rom_memory[3566] = 3'b100;
        rom_memory[3567] = 3'b100;
        rom_memory[3568] = 3'b100;
        rom_memory[3569] = 3'b100;
        rom_memory[3570] = 3'b100;
        rom_memory[3571] = 3'b100;
        rom_memory[3572] = 3'b100;
        rom_memory[3573] = 3'b100;
        rom_memory[3574] = 3'b100;
        rom_memory[3575] = 3'b110;
        rom_memory[3576] = 3'b110;
        rom_memory[3577] = 3'b100;
        rom_memory[3578] = 3'b100;
        rom_memory[3579] = 3'b100;
        rom_memory[3580] = 3'b100;
        rom_memory[3581] = 3'b100;
        rom_memory[3582] = 3'b100;
        rom_memory[3583] = 3'b100;
        rom_memory[3584] = 3'b110;
        rom_memory[3585] = 3'b100;
        rom_memory[3586] = 3'b100;
        rom_memory[3587] = 3'b110;
        rom_memory[3588] = 3'b100;
        rom_memory[3589] = 3'b100;
        rom_memory[3590] = 3'b110;
        rom_memory[3591] = 3'b110;
        rom_memory[3592] = 3'b100;
        rom_memory[3593] = 3'b110;
        rom_memory[3594] = 3'b110;
        rom_memory[3595] = 3'b110;
        rom_memory[3596] = 3'b110;
        rom_memory[3597] = 3'b110;
        rom_memory[3598] = 3'b110;
        rom_memory[3599] = 3'b110;
        rom_memory[3600] = 3'b110;
        rom_memory[3601] = 3'b110;
        rom_memory[3602] = 3'b110;
        rom_memory[3603] = 3'b110;
        rom_memory[3604] = 3'b110;
        rom_memory[3605] = 3'b110;
        rom_memory[3606] = 3'b110;
        rom_memory[3607] = 3'b110;
        rom_memory[3608] = 3'b110;
        rom_memory[3609] = 3'b110;
        rom_memory[3610] = 3'b110;
        rom_memory[3611] = 3'b110;
        rom_memory[3612] = 3'b110;
        rom_memory[3613] = 3'b110;
        rom_memory[3614] = 3'b110;
        rom_memory[3615] = 3'b110;
        rom_memory[3616] = 3'b110;
        rom_memory[3617] = 3'b110;
        rom_memory[3618] = 3'b110;
        rom_memory[3619] = 3'b110;
        rom_memory[3620] = 3'b110;
        rom_memory[3621] = 3'b110;
        rom_memory[3622] = 3'b110;
        rom_memory[3623] = 3'b110;
        rom_memory[3624] = 3'b110;
        rom_memory[3625] = 3'b110;
        rom_memory[3626] = 3'b110;
        rom_memory[3627] = 3'b110;
        rom_memory[3628] = 3'b110;
        rom_memory[3629] = 3'b110;
        rom_memory[3630] = 3'b110;
        rom_memory[3631] = 3'b110;
        rom_memory[3632] = 3'b110;
        rom_memory[3633] = 3'b110;
        rom_memory[3634] = 3'b110;
        rom_memory[3635] = 3'b110;
        rom_memory[3636] = 3'b110;
        rom_memory[3637] = 3'b110;
        rom_memory[3638] = 3'b110;
        rom_memory[3639] = 3'b110;
        rom_memory[3640] = 3'b110;
        rom_memory[3641] = 3'b110;
        rom_memory[3642] = 3'b110;
        rom_memory[3643] = 3'b110;
        rom_memory[3644] = 3'b110;
        rom_memory[3645] = 3'b110;
        rom_memory[3646] = 3'b110;
        rom_memory[3647] = 3'b110;
        rom_memory[3648] = 3'b110;
        rom_memory[3649] = 3'b110;
        rom_memory[3650] = 3'b110;
        rom_memory[3651] = 3'b110;
        rom_memory[3652] = 3'b110;
        rom_memory[3653] = 3'b110;
        rom_memory[3654] = 3'b110;
        rom_memory[3655] = 3'b110;
        rom_memory[3656] = 3'b110;
        rom_memory[3657] = 3'b110;
        rom_memory[3658] = 3'b110;
        rom_memory[3659] = 3'b110;
        rom_memory[3660] = 3'b110;
        rom_memory[3661] = 3'b110;
        rom_memory[3662] = 3'b110;
        rom_memory[3663] = 3'b110;
        rom_memory[3664] = 3'b110;
        rom_memory[3665] = 3'b110;
        rom_memory[3666] = 3'b110;
        rom_memory[3667] = 3'b110;
        rom_memory[3668] = 3'b110;
        rom_memory[3669] = 3'b110;
        rom_memory[3670] = 3'b110;
        rom_memory[3671] = 3'b110;
        rom_memory[3672] = 3'b110;
        rom_memory[3673] = 3'b110;
        rom_memory[3674] = 3'b110;
        rom_memory[3675] = 3'b110;
        rom_memory[3676] = 3'b110;
        rom_memory[3677] = 3'b110;
        rom_memory[3678] = 3'b110;
        rom_memory[3679] = 3'b110;
        rom_memory[3680] = 3'b110;
        rom_memory[3681] = 3'b110;
        rom_memory[3682] = 3'b110;
        rom_memory[3683] = 3'b110;
        rom_memory[3684] = 3'b110;
        rom_memory[3685] = 3'b110;
        rom_memory[3686] = 3'b110;
        rom_memory[3687] = 3'b110;
        rom_memory[3688] = 3'b110;
        rom_memory[3689] = 3'b110;
        rom_memory[3690] = 3'b110;
        rom_memory[3691] = 3'b110;
        rom_memory[3692] = 3'b110;
        rom_memory[3693] = 3'b110;
        rom_memory[3694] = 3'b110;
        rom_memory[3695] = 3'b110;
        rom_memory[3696] = 3'b110;
        rom_memory[3697] = 3'b110;
        rom_memory[3698] = 3'b110;
        rom_memory[3699] = 3'b110;
        rom_memory[3700] = 3'b110;
        rom_memory[3701] = 3'b110;
        rom_memory[3702] = 3'b110;
        rom_memory[3703] = 3'b110;
        rom_memory[3704] = 3'b110;
        rom_memory[3705] = 3'b110;
        rom_memory[3706] = 3'b110;
        rom_memory[3707] = 3'b110;
        rom_memory[3708] = 3'b110;
        rom_memory[3709] = 3'b110;
        rom_memory[3710] = 3'b110;
        rom_memory[3711] = 3'b110;
        rom_memory[3712] = 3'b110;
        rom_memory[3713] = 3'b110;
        rom_memory[3714] = 3'b110;
        rom_memory[3715] = 3'b110;
        rom_memory[3716] = 3'b110;
        rom_memory[3717] = 3'b110;
        rom_memory[3718] = 3'b110;
        rom_memory[3719] = 3'b110;
        rom_memory[3720] = 3'b110;
        rom_memory[3721] = 3'b110;
        rom_memory[3722] = 3'b110;
        rom_memory[3723] = 3'b110;
        rom_memory[3724] = 3'b110;
        rom_memory[3725] = 3'b110;
        rom_memory[3726] = 3'b110;
        rom_memory[3727] = 3'b110;
        rom_memory[3728] = 3'b110;
        rom_memory[3729] = 3'b110;
        rom_memory[3730] = 3'b110;
        rom_memory[3731] = 3'b110;
        rom_memory[3732] = 3'b110;
        rom_memory[3733] = 3'b110;
        rom_memory[3734] = 3'b110;
        rom_memory[3735] = 3'b110;
        rom_memory[3736] = 3'b110;
        rom_memory[3737] = 3'b110;
        rom_memory[3738] = 3'b110;
        rom_memory[3739] = 3'b110;
        rom_memory[3740] = 3'b110;
        rom_memory[3741] = 3'b110;
        rom_memory[3742] = 3'b110;
        rom_memory[3743] = 3'b110;
        rom_memory[3744] = 3'b110;
        rom_memory[3745] = 3'b110;
        rom_memory[3746] = 3'b110;
        rom_memory[3747] = 3'b110;
        rom_memory[3748] = 3'b110;
        rom_memory[3749] = 3'b110;
        rom_memory[3750] = 3'b110;
        rom_memory[3751] = 3'b110;
        rom_memory[3752] = 3'b110;
        rom_memory[3753] = 3'b110;
        rom_memory[3754] = 3'b110;
        rom_memory[3755] = 3'b110;
        rom_memory[3756] = 3'b110;
        rom_memory[3757] = 3'b110;
        rom_memory[3758] = 3'b110;
        rom_memory[3759] = 3'b110;
        rom_memory[3760] = 3'b110;
        rom_memory[3761] = 3'b110;
        rom_memory[3762] = 3'b110;
        rom_memory[3763] = 3'b110;
        rom_memory[3764] = 3'b110;
        rom_memory[3765] = 3'b110;
        rom_memory[3766] = 3'b110;
        rom_memory[3767] = 3'b110;
        rom_memory[3768] = 3'b110;
        rom_memory[3769] = 3'b100;
        rom_memory[3770] = 3'b110;
        rom_memory[3771] = 3'b100;
        rom_memory[3772] = 3'b110;
        rom_memory[3773] = 3'b110;
        rom_memory[3774] = 3'b110;
        rom_memory[3775] = 3'b110;
        rom_memory[3776] = 3'b110;
        rom_memory[3777] = 3'b100;
        rom_memory[3778] = 3'b100;
        rom_memory[3779] = 3'b100;
        rom_memory[3780] = 3'b100;
        rom_memory[3781] = 3'b100;
        rom_memory[3782] = 3'b100;
        rom_memory[3783] = 3'b100;
        rom_memory[3784] = 3'b100;
        rom_memory[3785] = 3'b100;
        rom_memory[3786] = 3'b100;
        rom_memory[3787] = 3'b110;
        rom_memory[3788] = 3'b100;
        rom_memory[3789] = 3'b110;
        rom_memory[3790] = 3'b100;
        rom_memory[3791] = 3'b110;
        rom_memory[3792] = 3'b110;
        rom_memory[3793] = 3'b100;
        rom_memory[3794] = 3'b100;
        rom_memory[3795] = 3'b100;
        rom_memory[3796] = 3'b100;
        rom_memory[3797] = 3'b100;
        rom_memory[3798] = 3'b110;
        rom_memory[3799] = 3'b110;
        rom_memory[3800] = 3'b110;
        rom_memory[3801] = 3'b110;
        rom_memory[3802] = 3'b100;
        rom_memory[3803] = 3'b100;
        rom_memory[3804] = 3'b100;
        rom_memory[3805] = 3'b100;
        rom_memory[3806] = 3'b100;
        rom_memory[3807] = 3'b100;
        rom_memory[3808] = 3'b100;
        rom_memory[3809] = 3'b100;
        rom_memory[3810] = 3'b100;
        rom_memory[3811] = 3'b100;
        rom_memory[3812] = 3'b100;
        rom_memory[3813] = 3'b100;
        rom_memory[3814] = 3'b100;
        rom_memory[3815] = 3'b110;
        rom_memory[3816] = 3'b110;
        rom_memory[3817] = 3'b100;
        rom_memory[3818] = 3'b100;
        rom_memory[3819] = 3'b110;
        rom_memory[3820] = 3'b100;
        rom_memory[3821] = 3'b100;
        rom_memory[3822] = 3'b100;
        rom_memory[3823] = 3'b100;
        rom_memory[3824] = 3'b110;
        rom_memory[3825] = 3'b110;
        rom_memory[3826] = 3'b110;
        rom_memory[3827] = 3'b110;
        rom_memory[3828] = 3'b110;
        rom_memory[3829] = 3'b110;
        rom_memory[3830] = 3'b100;
        rom_memory[3831] = 3'b110;
        rom_memory[3832] = 3'b110;
        rom_memory[3833] = 3'b110;
        rom_memory[3834] = 3'b110;
        rom_memory[3835] = 3'b110;
        rom_memory[3836] = 3'b110;
        rom_memory[3837] = 3'b110;
        rom_memory[3838] = 3'b110;
        rom_memory[3839] = 3'b110;
        rom_memory[3840] = 3'b110;
        rom_memory[3841] = 3'b110;
        rom_memory[3842] = 3'b110;
        rom_memory[3843] = 3'b110;
        rom_memory[3844] = 3'b110;
        rom_memory[3845] = 3'b110;
        rom_memory[3846] = 3'b110;
        rom_memory[3847] = 3'b110;
        rom_memory[3848] = 3'b110;
        rom_memory[3849] = 3'b110;
        rom_memory[3850] = 3'b110;
        rom_memory[3851] = 3'b110;
        rom_memory[3852] = 3'b110;
        rom_memory[3853] = 3'b110;
        rom_memory[3854] = 3'b110;
        rom_memory[3855] = 3'b110;
        rom_memory[3856] = 3'b110;
        rom_memory[3857] = 3'b110;
        rom_memory[3858] = 3'b110;
        rom_memory[3859] = 3'b110;
        rom_memory[3860] = 3'b110;
        rom_memory[3861] = 3'b110;
        rom_memory[3862] = 3'b110;
        rom_memory[3863] = 3'b110;
        rom_memory[3864] = 3'b110;
        rom_memory[3865] = 3'b110;
        rom_memory[3866] = 3'b110;
        rom_memory[3867] = 3'b110;
        rom_memory[3868] = 3'b110;
        rom_memory[3869] = 3'b110;
        rom_memory[3870] = 3'b110;
        rom_memory[3871] = 3'b110;
        rom_memory[3872] = 3'b110;
        rom_memory[3873] = 3'b110;
        rom_memory[3874] = 3'b110;
        rom_memory[3875] = 3'b110;
        rom_memory[3876] = 3'b110;
        rom_memory[3877] = 3'b110;
        rom_memory[3878] = 3'b110;
        rom_memory[3879] = 3'b110;
        rom_memory[3880] = 3'b110;
        rom_memory[3881] = 3'b110;
        rom_memory[3882] = 3'b110;
        rom_memory[3883] = 3'b110;
        rom_memory[3884] = 3'b110;
        rom_memory[3885] = 3'b110;
        rom_memory[3886] = 3'b110;
        rom_memory[3887] = 3'b110;
        rom_memory[3888] = 3'b110;
        rom_memory[3889] = 3'b110;
        rom_memory[3890] = 3'b110;
        rom_memory[3891] = 3'b110;
        rom_memory[3892] = 3'b110;
        rom_memory[3893] = 3'b110;
        rom_memory[3894] = 3'b110;
        rom_memory[3895] = 3'b110;
        rom_memory[3896] = 3'b110;
        rom_memory[3897] = 3'b110;
        rom_memory[3898] = 3'b110;
        rom_memory[3899] = 3'b110;
        rom_memory[3900] = 3'b110;
        rom_memory[3901] = 3'b110;
        rom_memory[3902] = 3'b110;
        rom_memory[3903] = 3'b110;
        rom_memory[3904] = 3'b110;
        rom_memory[3905] = 3'b110;
        rom_memory[3906] = 3'b110;
        rom_memory[3907] = 3'b110;
        rom_memory[3908] = 3'b110;
        rom_memory[3909] = 3'b110;
        rom_memory[3910] = 3'b110;
        rom_memory[3911] = 3'b110;
        rom_memory[3912] = 3'b110;
        rom_memory[3913] = 3'b110;
        rom_memory[3914] = 3'b110;
        rom_memory[3915] = 3'b110;
        rom_memory[3916] = 3'b110;
        rom_memory[3917] = 3'b110;
        rom_memory[3918] = 3'b110;
        rom_memory[3919] = 3'b110;
        rom_memory[3920] = 3'b110;
        rom_memory[3921] = 3'b110;
        rom_memory[3922] = 3'b110;
        rom_memory[3923] = 3'b110;
        rom_memory[3924] = 3'b110;
        rom_memory[3925] = 3'b110;
        rom_memory[3926] = 3'b110;
        rom_memory[3927] = 3'b110;
        rom_memory[3928] = 3'b110;
        rom_memory[3929] = 3'b110;
        rom_memory[3930] = 3'b110;
        rom_memory[3931] = 3'b110;
        rom_memory[3932] = 3'b110;
        rom_memory[3933] = 3'b110;
        rom_memory[3934] = 3'b110;
        rom_memory[3935] = 3'b110;
        rom_memory[3936] = 3'b110;
        rom_memory[3937] = 3'b110;
        rom_memory[3938] = 3'b110;
        rom_memory[3939] = 3'b110;
        rom_memory[3940] = 3'b110;
        rom_memory[3941] = 3'b110;
        rom_memory[3942] = 3'b110;
        rom_memory[3943] = 3'b110;
        rom_memory[3944] = 3'b110;
        rom_memory[3945] = 3'b110;
        rom_memory[3946] = 3'b110;
        rom_memory[3947] = 3'b110;
        rom_memory[3948] = 3'b110;
        rom_memory[3949] = 3'b110;
        rom_memory[3950] = 3'b110;
        rom_memory[3951] = 3'b110;
        rom_memory[3952] = 3'b110;
        rom_memory[3953] = 3'b110;
        rom_memory[3954] = 3'b110;
        rom_memory[3955] = 3'b110;
        rom_memory[3956] = 3'b110;
        rom_memory[3957] = 3'b110;
        rom_memory[3958] = 3'b110;
        rom_memory[3959] = 3'b110;
        rom_memory[3960] = 3'b110;
        rom_memory[3961] = 3'b110;
        rom_memory[3962] = 3'b110;
        rom_memory[3963] = 3'b110;
        rom_memory[3964] = 3'b110;
        rom_memory[3965] = 3'b110;
        rom_memory[3966] = 3'b110;
        rom_memory[3967] = 3'b110;
        rom_memory[3968] = 3'b110;
        rom_memory[3969] = 3'b110;
        rom_memory[3970] = 3'b110;
        rom_memory[3971] = 3'b110;
        rom_memory[3972] = 3'b110;
        rom_memory[3973] = 3'b110;
        rom_memory[3974] = 3'b110;
        rom_memory[3975] = 3'b110;
        rom_memory[3976] = 3'b110;
        rom_memory[3977] = 3'b110;
        rom_memory[3978] = 3'b110;
        rom_memory[3979] = 3'b110;
        rom_memory[3980] = 3'b110;
        rom_memory[3981] = 3'b110;
        rom_memory[3982] = 3'b110;
        rom_memory[3983] = 3'b110;
        rom_memory[3984] = 3'b110;
        rom_memory[3985] = 3'b110;
        rom_memory[3986] = 3'b110;
        rom_memory[3987] = 3'b110;
        rom_memory[3988] = 3'b110;
        rom_memory[3989] = 3'b110;
        rom_memory[3990] = 3'b110;
        rom_memory[3991] = 3'b110;
        rom_memory[3992] = 3'b110;
        rom_memory[3993] = 3'b110;
        rom_memory[3994] = 3'b110;
        rom_memory[3995] = 3'b110;
        rom_memory[3996] = 3'b110;
        rom_memory[3997] = 3'b110;
        rom_memory[3998] = 3'b110;
        rom_memory[3999] = 3'b110;
        rom_memory[4000] = 3'b110;
        rom_memory[4001] = 3'b110;
        rom_memory[4002] = 3'b110;
        rom_memory[4003] = 3'b110;
        rom_memory[4004] = 3'b110;
        rom_memory[4005] = 3'b110;
        rom_memory[4006] = 3'b110;
        rom_memory[4007] = 3'b110;
        rom_memory[4008] = 3'b110;
        rom_memory[4009] = 3'b110;
        rom_memory[4010] = 3'b110;
        rom_memory[4011] = 3'b110;
        rom_memory[4012] = 3'b110;
        rom_memory[4013] = 3'b110;
        rom_memory[4014] = 3'b110;
        rom_memory[4015] = 3'b110;
        rom_memory[4016] = 3'b100;
        rom_memory[4017] = 3'b110;
        rom_memory[4018] = 3'b110;
        rom_memory[4019] = 3'b100;
        rom_memory[4020] = 3'b100;
        rom_memory[4021] = 3'b110;
        rom_memory[4022] = 3'b100;
        rom_memory[4023] = 3'b110;
        rom_memory[4024] = 3'b110;
        rom_memory[4025] = 3'b110;
        rom_memory[4026] = 3'b110;
        rom_memory[4027] = 3'b110;
        rom_memory[4028] = 3'b110;
        rom_memory[4029] = 3'b110;
        rom_memory[4030] = 3'b110;
        rom_memory[4031] = 3'b110;
        rom_memory[4032] = 3'b110;
        rom_memory[4033] = 3'b110;
        rom_memory[4034] = 3'b100;
        rom_memory[4035] = 3'b110;
        rom_memory[4036] = 3'b110;
        rom_memory[4037] = 3'b110;
        rom_memory[4038] = 3'b110;
        rom_memory[4039] = 3'b110;
        rom_memory[4040] = 3'b110;
        rom_memory[4041] = 3'b110;
        rom_memory[4042] = 3'b110;
        rom_memory[4043] = 3'b110;
        rom_memory[4044] = 3'b110;
        rom_memory[4045] = 3'b110;
        rom_memory[4046] = 3'b110;
        rom_memory[4047] = 3'b110;
        rom_memory[4048] = 3'b110;
        rom_memory[4049] = 3'b110;
        rom_memory[4050] = 3'b100;
        rom_memory[4051] = 3'b110;
        rom_memory[4052] = 3'b110;
        rom_memory[4053] = 3'b100;
        rom_memory[4054] = 3'b100;
        rom_memory[4055] = 3'b110;
        rom_memory[4056] = 3'b110;
        rom_memory[4057] = 3'b110;
        rom_memory[4058] = 3'b110;
        rom_memory[4059] = 3'b110;
        rom_memory[4060] = 3'b110;
        rom_memory[4061] = 3'b110;
        rom_memory[4062] = 3'b100;
        rom_memory[4063] = 3'b110;
        rom_memory[4064] = 3'b110;
        rom_memory[4065] = 3'b110;
        rom_memory[4066] = 3'b110;
        rom_memory[4067] = 3'b110;
        rom_memory[4068] = 3'b110;
        rom_memory[4069] = 3'b110;
        rom_memory[4070] = 3'b110;
        rom_memory[4071] = 3'b110;
        rom_memory[4072] = 3'b110;
        rom_memory[4073] = 3'b110;
        rom_memory[4074] = 3'b110;
        rom_memory[4075] = 3'b110;
        rom_memory[4076] = 3'b110;
        rom_memory[4077] = 3'b110;
        rom_memory[4078] = 3'b110;
        rom_memory[4079] = 3'b110;
        rom_memory[4080] = 3'b110;
        rom_memory[4081] = 3'b110;
        rom_memory[4082] = 3'b110;
        rom_memory[4083] = 3'b110;
        rom_memory[4084] = 3'b110;
        rom_memory[4085] = 3'b110;
        rom_memory[4086] = 3'b110;
        rom_memory[4087] = 3'b110;
        rom_memory[4088] = 3'b110;
        rom_memory[4089] = 3'b110;
        rom_memory[4090] = 3'b110;
        rom_memory[4091] = 3'b110;
        rom_memory[4092] = 3'b110;
        rom_memory[4093] = 3'b110;
        rom_memory[4094] = 3'b110;
        rom_memory[4095] = 3'b110;
        rom_memory[4096] = 3'b110;
        rom_memory[4097] = 3'b110;
        rom_memory[4098] = 3'b110;
        rom_memory[4099] = 3'b110;
        rom_memory[4100] = 3'b110;
        rom_memory[4101] = 3'b110;
        rom_memory[4102] = 3'b110;
        rom_memory[4103] = 3'b110;
        rom_memory[4104] = 3'b110;
        rom_memory[4105] = 3'b110;
        rom_memory[4106] = 3'b110;
        rom_memory[4107] = 3'b110;
        rom_memory[4108] = 3'b110;
        rom_memory[4109] = 3'b110;
        rom_memory[4110] = 3'b110;
        rom_memory[4111] = 3'b110;
        rom_memory[4112] = 3'b110;
        rom_memory[4113] = 3'b110;
        rom_memory[4114] = 3'b110;
        rom_memory[4115] = 3'b110;
        rom_memory[4116] = 3'b110;
        rom_memory[4117] = 3'b110;
        rom_memory[4118] = 3'b110;
        rom_memory[4119] = 3'b110;
        rom_memory[4120] = 3'b110;
        rom_memory[4121] = 3'b110;
        rom_memory[4122] = 3'b110;
        rom_memory[4123] = 3'b110;
        rom_memory[4124] = 3'b110;
        rom_memory[4125] = 3'b110;
        rom_memory[4126] = 3'b110;
        rom_memory[4127] = 3'b110;
        rom_memory[4128] = 3'b110;
        rom_memory[4129] = 3'b110;
        rom_memory[4130] = 3'b110;
        rom_memory[4131] = 3'b110;
        rom_memory[4132] = 3'b110;
        rom_memory[4133] = 3'b110;
        rom_memory[4134] = 3'b110;
        rom_memory[4135] = 3'b110;
        rom_memory[4136] = 3'b110;
        rom_memory[4137] = 3'b110;
        rom_memory[4138] = 3'b110;
        rom_memory[4139] = 3'b110;
        rom_memory[4140] = 3'b110;
        rom_memory[4141] = 3'b110;
        rom_memory[4142] = 3'b110;
        rom_memory[4143] = 3'b110;
        rom_memory[4144] = 3'b110;
        rom_memory[4145] = 3'b110;
        rom_memory[4146] = 3'b110;
        rom_memory[4147] = 3'b110;
        rom_memory[4148] = 3'b110;
        rom_memory[4149] = 3'b110;
        rom_memory[4150] = 3'b110;
        rom_memory[4151] = 3'b110;
        rom_memory[4152] = 3'b110;
        rom_memory[4153] = 3'b110;
        rom_memory[4154] = 3'b110;
        rom_memory[4155] = 3'b110;
        rom_memory[4156] = 3'b110;
        rom_memory[4157] = 3'b110;
        rom_memory[4158] = 3'b110;
        rom_memory[4159] = 3'b110;
        rom_memory[4160] = 3'b110;
        rom_memory[4161] = 3'b110;
        rom_memory[4162] = 3'b110;
        rom_memory[4163] = 3'b110;
        rom_memory[4164] = 3'b110;
        rom_memory[4165] = 3'b110;
        rom_memory[4166] = 3'b110;
        rom_memory[4167] = 3'b110;
        rom_memory[4168] = 3'b110;
        rom_memory[4169] = 3'b110;
        rom_memory[4170] = 3'b110;
        rom_memory[4171] = 3'b110;
        rom_memory[4172] = 3'b110;
        rom_memory[4173] = 3'b110;
        rom_memory[4174] = 3'b110;
        rom_memory[4175] = 3'b110;
        rom_memory[4176] = 3'b110;
        rom_memory[4177] = 3'b110;
        rom_memory[4178] = 3'b110;
        rom_memory[4179] = 3'b110;
        rom_memory[4180] = 3'b110;
        rom_memory[4181] = 3'b110;
        rom_memory[4182] = 3'b110;
        rom_memory[4183] = 3'b110;
        rom_memory[4184] = 3'b110;
        rom_memory[4185] = 3'b110;
        rom_memory[4186] = 3'b110;
        rom_memory[4187] = 3'b110;
        rom_memory[4188] = 3'b110;
        rom_memory[4189] = 3'b110;
        rom_memory[4190] = 3'b110;
        rom_memory[4191] = 3'b110;
        rom_memory[4192] = 3'b110;
        rom_memory[4193] = 3'b110;
        rom_memory[4194] = 3'b110;
        rom_memory[4195] = 3'b110;
        rom_memory[4196] = 3'b110;
        rom_memory[4197] = 3'b110;
        rom_memory[4198] = 3'b110;
        rom_memory[4199] = 3'b110;
        rom_memory[4200] = 3'b110;
        rom_memory[4201] = 3'b110;
        rom_memory[4202] = 3'b110;
        rom_memory[4203] = 3'b110;
        rom_memory[4204] = 3'b110;
        rom_memory[4205] = 3'b110;
        rom_memory[4206] = 3'b110;
        rom_memory[4207] = 3'b110;
        rom_memory[4208] = 3'b110;
        rom_memory[4209] = 3'b110;
        rom_memory[4210] = 3'b110;
        rom_memory[4211] = 3'b110;
        rom_memory[4212] = 3'b110;
        rom_memory[4213] = 3'b110;
        rom_memory[4214] = 3'b110;
        rom_memory[4215] = 3'b110;
        rom_memory[4216] = 3'b110;
        rom_memory[4217] = 3'b110;
        rom_memory[4218] = 3'b110;
        rom_memory[4219] = 3'b110;
        rom_memory[4220] = 3'b110;
        rom_memory[4221] = 3'b110;
        rom_memory[4222] = 3'b110;
        rom_memory[4223] = 3'b110;
        rom_memory[4224] = 3'b110;
        rom_memory[4225] = 3'b110;
        rom_memory[4226] = 3'b110;
        rom_memory[4227] = 3'b110;
        rom_memory[4228] = 3'b110;
        rom_memory[4229] = 3'b110;
        rom_memory[4230] = 3'b110;
        rom_memory[4231] = 3'b110;
        rom_memory[4232] = 3'b110;
        rom_memory[4233] = 3'b110;
        rom_memory[4234] = 3'b110;
        rom_memory[4235] = 3'b110;
        rom_memory[4236] = 3'b110;
        rom_memory[4237] = 3'b110;
        rom_memory[4238] = 3'b110;
        rom_memory[4239] = 3'b110;
        rom_memory[4240] = 3'b110;
        rom_memory[4241] = 3'b110;
        rom_memory[4242] = 3'b110;
        rom_memory[4243] = 3'b110;
        rom_memory[4244] = 3'b110;
        rom_memory[4245] = 3'b110;
        rom_memory[4246] = 3'b110;
        rom_memory[4247] = 3'b110;
        rom_memory[4248] = 3'b110;
        rom_memory[4249] = 3'b110;
        rom_memory[4250] = 3'b110;
        rom_memory[4251] = 3'b110;
        rom_memory[4252] = 3'b110;
        rom_memory[4253] = 3'b110;
        rom_memory[4254] = 3'b110;
        rom_memory[4255] = 3'b110;
        rom_memory[4256] = 3'b110;
        rom_memory[4257] = 3'b110;
        rom_memory[4258] = 3'b110;
        rom_memory[4259] = 3'b110;
        rom_memory[4260] = 3'b110;
        rom_memory[4261] = 3'b110;
        rom_memory[4262] = 3'b110;
        rom_memory[4263] = 3'b110;
        rom_memory[4264] = 3'b110;
        rom_memory[4265] = 3'b110;
        rom_memory[4266] = 3'b110;
        rom_memory[4267] = 3'b110;
        rom_memory[4268] = 3'b110;
        rom_memory[4269] = 3'b110;
        rom_memory[4270] = 3'b110;
        rom_memory[4271] = 3'b110;
        rom_memory[4272] = 3'b110;
        rom_memory[4273] = 3'b110;
        rom_memory[4274] = 3'b110;
        rom_memory[4275] = 3'b110;
        rom_memory[4276] = 3'b110;
        rom_memory[4277] = 3'b110;
        rom_memory[4278] = 3'b110;
        rom_memory[4279] = 3'b110;
        rom_memory[4280] = 3'b110;
        rom_memory[4281] = 3'b110;
        rom_memory[4282] = 3'b110;
        rom_memory[4283] = 3'b110;
        rom_memory[4284] = 3'b110;
        rom_memory[4285] = 3'b110;
        rom_memory[4286] = 3'b110;
        rom_memory[4287] = 3'b110;
        rom_memory[4288] = 3'b110;
        rom_memory[4289] = 3'b110;
        rom_memory[4290] = 3'b110;
        rom_memory[4291] = 3'b110;
        rom_memory[4292] = 3'b110;
        rom_memory[4293] = 3'b110;
        rom_memory[4294] = 3'b110;
        rom_memory[4295] = 3'b110;
        rom_memory[4296] = 3'b110;
        rom_memory[4297] = 3'b110;
        rom_memory[4298] = 3'b110;
        rom_memory[4299] = 3'b110;
        rom_memory[4300] = 3'b110;
        rom_memory[4301] = 3'b110;
        rom_memory[4302] = 3'b110;
        rom_memory[4303] = 3'b110;
        rom_memory[4304] = 3'b110;
        rom_memory[4305] = 3'b110;
        rom_memory[4306] = 3'b110;
        rom_memory[4307] = 3'b110;
        rom_memory[4308] = 3'b110;
        rom_memory[4309] = 3'b110;
        rom_memory[4310] = 3'b110;
        rom_memory[4311] = 3'b110;
        rom_memory[4312] = 3'b110;
        rom_memory[4313] = 3'b110;
        rom_memory[4314] = 3'b110;
        rom_memory[4315] = 3'b110;
        rom_memory[4316] = 3'b110;
        rom_memory[4317] = 3'b110;
        rom_memory[4318] = 3'b110;
        rom_memory[4319] = 3'b110;
        rom_memory[4320] = 3'b110;
        rom_memory[4321] = 3'b110;
        rom_memory[4322] = 3'b110;
        rom_memory[4323] = 3'b110;
        rom_memory[4324] = 3'b110;
        rom_memory[4325] = 3'b110;
        rom_memory[4326] = 3'b110;
        rom_memory[4327] = 3'b110;
        rom_memory[4328] = 3'b110;
        rom_memory[4329] = 3'b110;
        rom_memory[4330] = 3'b110;
        rom_memory[4331] = 3'b110;
        rom_memory[4332] = 3'b110;
        rom_memory[4333] = 3'b110;
        rom_memory[4334] = 3'b110;
        rom_memory[4335] = 3'b110;
        rom_memory[4336] = 3'b110;
        rom_memory[4337] = 3'b110;
        rom_memory[4338] = 3'b110;
        rom_memory[4339] = 3'b110;
        rom_memory[4340] = 3'b110;
        rom_memory[4341] = 3'b110;
        rom_memory[4342] = 3'b110;
        rom_memory[4343] = 3'b110;
        rom_memory[4344] = 3'b110;
        rom_memory[4345] = 3'b110;
        rom_memory[4346] = 3'b110;
        rom_memory[4347] = 3'b110;
        rom_memory[4348] = 3'b110;
        rom_memory[4349] = 3'b110;
        rom_memory[4350] = 3'b110;
        rom_memory[4351] = 3'b110;
        rom_memory[4352] = 3'b110;
        rom_memory[4353] = 3'b110;
        rom_memory[4354] = 3'b110;
        rom_memory[4355] = 3'b110;
        rom_memory[4356] = 3'b110;
        rom_memory[4357] = 3'b110;
        rom_memory[4358] = 3'b110;
        rom_memory[4359] = 3'b110;
        rom_memory[4360] = 3'b110;
        rom_memory[4361] = 3'b110;
        rom_memory[4362] = 3'b110;
        rom_memory[4363] = 3'b110;
        rom_memory[4364] = 3'b110;
        rom_memory[4365] = 3'b110;
        rom_memory[4366] = 3'b110;
        rom_memory[4367] = 3'b110;
        rom_memory[4368] = 3'b110;
        rom_memory[4369] = 3'b110;
        rom_memory[4370] = 3'b110;
        rom_memory[4371] = 3'b110;
        rom_memory[4372] = 3'b110;
        rom_memory[4373] = 3'b110;
        rom_memory[4374] = 3'b110;
        rom_memory[4375] = 3'b110;
        rom_memory[4376] = 3'b110;
        rom_memory[4377] = 3'b110;
        rom_memory[4378] = 3'b110;
        rom_memory[4379] = 3'b110;
        rom_memory[4380] = 3'b110;
        rom_memory[4381] = 3'b110;
        rom_memory[4382] = 3'b110;
        rom_memory[4383] = 3'b110;
        rom_memory[4384] = 3'b110;
        rom_memory[4385] = 3'b110;
        rom_memory[4386] = 3'b110;
        rom_memory[4387] = 3'b110;
        rom_memory[4388] = 3'b110;
        rom_memory[4389] = 3'b110;
        rom_memory[4390] = 3'b110;
        rom_memory[4391] = 3'b110;
        rom_memory[4392] = 3'b110;
        rom_memory[4393] = 3'b110;
        rom_memory[4394] = 3'b110;
        rom_memory[4395] = 3'b110;
        rom_memory[4396] = 3'b110;
        rom_memory[4397] = 3'b110;
        rom_memory[4398] = 3'b110;
        rom_memory[4399] = 3'b110;
        rom_memory[4400] = 3'b110;
        rom_memory[4401] = 3'b110;
        rom_memory[4402] = 3'b110;
        rom_memory[4403] = 3'b110;
        rom_memory[4404] = 3'b110;
        rom_memory[4405] = 3'b110;
        rom_memory[4406] = 3'b110;
        rom_memory[4407] = 3'b110;
        rom_memory[4408] = 3'b110;
        rom_memory[4409] = 3'b110;
        rom_memory[4410] = 3'b110;
        rom_memory[4411] = 3'b110;
        rom_memory[4412] = 3'b110;
        rom_memory[4413] = 3'b110;
        rom_memory[4414] = 3'b110;
        rom_memory[4415] = 3'b110;
        rom_memory[4416] = 3'b110;
        rom_memory[4417] = 3'b110;
        rom_memory[4418] = 3'b110;
        rom_memory[4419] = 3'b110;
        rom_memory[4420] = 3'b110;
        rom_memory[4421] = 3'b110;
        rom_memory[4422] = 3'b110;
        rom_memory[4423] = 3'b110;
        rom_memory[4424] = 3'b110;
        rom_memory[4425] = 3'b110;
        rom_memory[4426] = 3'b110;
        rom_memory[4427] = 3'b110;
        rom_memory[4428] = 3'b110;
        rom_memory[4429] = 3'b110;
        rom_memory[4430] = 3'b110;
        rom_memory[4431] = 3'b110;
        rom_memory[4432] = 3'b110;
        rom_memory[4433] = 3'b110;
        rom_memory[4434] = 3'b110;
        rom_memory[4435] = 3'b110;
        rom_memory[4436] = 3'b110;
        rom_memory[4437] = 3'b110;
        rom_memory[4438] = 3'b110;
        rom_memory[4439] = 3'b110;
        rom_memory[4440] = 3'b110;
        rom_memory[4441] = 3'b110;
        rom_memory[4442] = 3'b110;
        rom_memory[4443] = 3'b110;
        rom_memory[4444] = 3'b110;
        rom_memory[4445] = 3'b110;
        rom_memory[4446] = 3'b110;
        rom_memory[4447] = 3'b110;
        rom_memory[4448] = 3'b110;
        rom_memory[4449] = 3'b110;
        rom_memory[4450] = 3'b110;
        rom_memory[4451] = 3'b110;
        rom_memory[4452] = 3'b110;
        rom_memory[4453] = 3'b110;
        rom_memory[4454] = 3'b110;
        rom_memory[4455] = 3'b110;
        rom_memory[4456] = 3'b110;
        rom_memory[4457] = 3'b110;
        rom_memory[4458] = 3'b110;
        rom_memory[4459] = 3'b110;
        rom_memory[4460] = 3'b110;
        rom_memory[4461] = 3'b110;
        rom_memory[4462] = 3'b110;
        rom_memory[4463] = 3'b110;
        rom_memory[4464] = 3'b110;
        rom_memory[4465] = 3'b110;
        rom_memory[4466] = 3'b110;
        rom_memory[4467] = 3'b110;
        rom_memory[4468] = 3'b110;
        rom_memory[4469] = 3'b110;
        rom_memory[4470] = 3'b110;
        rom_memory[4471] = 3'b110;
        rom_memory[4472] = 3'b110;
        rom_memory[4473] = 3'b110;
        rom_memory[4474] = 3'b110;
        rom_memory[4475] = 3'b110;
        rom_memory[4476] = 3'b110;
        rom_memory[4477] = 3'b110;
        rom_memory[4478] = 3'b110;
        rom_memory[4479] = 3'b110;
        rom_memory[4480] = 3'b110;
        rom_memory[4481] = 3'b110;
        rom_memory[4482] = 3'b110;
        rom_memory[4483] = 3'b110;
        rom_memory[4484] = 3'b110;
        rom_memory[4485] = 3'b110;
        rom_memory[4486] = 3'b110;
        rom_memory[4487] = 3'b110;
        rom_memory[4488] = 3'b110;
        rom_memory[4489] = 3'b110;
        rom_memory[4490] = 3'b110;
        rom_memory[4491] = 3'b110;
        rom_memory[4492] = 3'b110;
        rom_memory[4493] = 3'b110;
        rom_memory[4494] = 3'b110;
        rom_memory[4495] = 3'b110;
        rom_memory[4496] = 3'b110;
        rom_memory[4497] = 3'b110;
        rom_memory[4498] = 3'b110;
        rom_memory[4499] = 3'b110;
        rom_memory[4500] = 3'b110;
        rom_memory[4501] = 3'b110;
        rom_memory[4502] = 3'b110;
        rom_memory[4503] = 3'b110;
        rom_memory[4504] = 3'b110;
        rom_memory[4505] = 3'b110;
        rom_memory[4506] = 3'b110;
        rom_memory[4507] = 3'b110;
        rom_memory[4508] = 3'b110;
        rom_memory[4509] = 3'b110;
        rom_memory[4510] = 3'b110;
        rom_memory[4511] = 3'b110;
        rom_memory[4512] = 3'b110;
        rom_memory[4513] = 3'b110;
        rom_memory[4514] = 3'b110;
        rom_memory[4515] = 3'b110;
        rom_memory[4516] = 3'b110;
        rom_memory[4517] = 3'b110;
        rom_memory[4518] = 3'b110;
        rom_memory[4519] = 3'b110;
        rom_memory[4520] = 3'b110;
        rom_memory[4521] = 3'b110;
        rom_memory[4522] = 3'b110;
        rom_memory[4523] = 3'b110;
        rom_memory[4524] = 3'b110;
        rom_memory[4525] = 3'b110;
        rom_memory[4526] = 3'b110;
        rom_memory[4527] = 3'b110;
        rom_memory[4528] = 3'b110;
        rom_memory[4529] = 3'b110;
        rom_memory[4530] = 3'b110;
        rom_memory[4531] = 3'b110;
        rom_memory[4532] = 3'b110;
        rom_memory[4533] = 3'b110;
        rom_memory[4534] = 3'b110;
        rom_memory[4535] = 3'b110;
        rom_memory[4536] = 3'b110;
        rom_memory[4537] = 3'b110;
        rom_memory[4538] = 3'b110;
        rom_memory[4539] = 3'b110;
        rom_memory[4540] = 3'b110;
        rom_memory[4541] = 3'b110;
        rom_memory[4542] = 3'b110;
        rom_memory[4543] = 3'b110;
        rom_memory[4544] = 3'b110;
        rom_memory[4545] = 3'b110;
        rom_memory[4546] = 3'b110;
        rom_memory[4547] = 3'b110;
        rom_memory[4548] = 3'b110;
        rom_memory[4549] = 3'b110;
        rom_memory[4550] = 3'b110;
        rom_memory[4551] = 3'b110;
        rom_memory[4552] = 3'b110;
        rom_memory[4553] = 3'b110;
        rom_memory[4554] = 3'b110;
        rom_memory[4555] = 3'b110;
        rom_memory[4556] = 3'b110;
        rom_memory[4557] = 3'b110;
        rom_memory[4558] = 3'b110;
        rom_memory[4559] = 3'b110;
        rom_memory[4560] = 3'b110;
        rom_memory[4561] = 3'b110;
        rom_memory[4562] = 3'b110;
        rom_memory[4563] = 3'b110;
        rom_memory[4564] = 3'b110;
        rom_memory[4565] = 3'b110;
        rom_memory[4566] = 3'b110;
        rom_memory[4567] = 3'b110;
        rom_memory[4568] = 3'b110;
        rom_memory[4569] = 3'b110;
        rom_memory[4570] = 3'b110;
        rom_memory[4571] = 3'b110;
        rom_memory[4572] = 3'b110;
        rom_memory[4573] = 3'b110;
        rom_memory[4574] = 3'b110;
        rom_memory[4575] = 3'b110;
        rom_memory[4576] = 3'b110;
        rom_memory[4577] = 3'b110;
        rom_memory[4578] = 3'b110;
        rom_memory[4579] = 3'b110;
        rom_memory[4580] = 3'b111;
        rom_memory[4581] = 3'b111;
        rom_memory[4582] = 3'b111;
        rom_memory[4583] = 3'b111;
        rom_memory[4584] = 3'b111;
        rom_memory[4585] = 3'b111;
        rom_memory[4586] = 3'b111;
        rom_memory[4587] = 3'b111;
        rom_memory[4588] = 3'b111;
        rom_memory[4589] = 3'b111;
        rom_memory[4590] = 3'b110;
        rom_memory[4591] = 3'b110;
        rom_memory[4592] = 3'b110;
        rom_memory[4593] = 3'b110;
        rom_memory[4594] = 3'b110;
        rom_memory[4595] = 3'b110;
        rom_memory[4596] = 3'b110;
        rom_memory[4597] = 3'b110;
        rom_memory[4598] = 3'b110;
        rom_memory[4599] = 3'b110;
        rom_memory[4600] = 3'b110;
        rom_memory[4601] = 3'b110;
        rom_memory[4602] = 3'b110;
        rom_memory[4603] = 3'b110;
        rom_memory[4604] = 3'b110;
        rom_memory[4605] = 3'b110;
        rom_memory[4606] = 3'b110;
        rom_memory[4607] = 3'b110;
        rom_memory[4608] = 3'b110;
        rom_memory[4609] = 3'b110;
        rom_memory[4610] = 3'b110;
        rom_memory[4611] = 3'b110;
        rom_memory[4612] = 3'b110;
        rom_memory[4613] = 3'b110;
        rom_memory[4614] = 3'b110;
        rom_memory[4615] = 3'b110;
        rom_memory[4616] = 3'b110;
        rom_memory[4617] = 3'b110;
        rom_memory[4618] = 3'b110;
        rom_memory[4619] = 3'b110;
        rom_memory[4620] = 3'b110;
        rom_memory[4621] = 3'b111;
        rom_memory[4622] = 3'b111;
        rom_memory[4623] = 3'b111;
        rom_memory[4624] = 3'b111;
        rom_memory[4625] = 3'b111;
        rom_memory[4626] = 3'b111;
        rom_memory[4627] = 3'b111;
        rom_memory[4628] = 3'b111;
        rom_memory[4629] = 3'b111;
        rom_memory[4630] = 3'b111;
        rom_memory[4631] = 3'b111;
        rom_memory[4632] = 3'b111;
        rom_memory[4633] = 3'b110;
        rom_memory[4634] = 3'b110;
        rom_memory[4635] = 3'b110;
        rom_memory[4636] = 3'b110;
        rom_memory[4637] = 3'b110;
        rom_memory[4638] = 3'b110;
        rom_memory[4639] = 3'b110;
        rom_memory[4640] = 3'b110;
        rom_memory[4641] = 3'b110;
        rom_memory[4642] = 3'b110;
        rom_memory[4643] = 3'b110;
        rom_memory[4644] = 3'b110;
        rom_memory[4645] = 3'b110;
        rom_memory[4646] = 3'b110;
        rom_memory[4647] = 3'b110;
        rom_memory[4648] = 3'b110;
        rom_memory[4649] = 3'b110;
        rom_memory[4650] = 3'b110;
        rom_memory[4651] = 3'b110;
        rom_memory[4652] = 3'b110;
        rom_memory[4653] = 3'b110;
        rom_memory[4654] = 3'b110;
        rom_memory[4655] = 3'b110;
        rom_memory[4656] = 3'b110;
        rom_memory[4657] = 3'b110;
        rom_memory[4658] = 3'b110;
        rom_memory[4659] = 3'b110;
        rom_memory[4660] = 3'b110;
        rom_memory[4661] = 3'b110;
        rom_memory[4662] = 3'b110;
        rom_memory[4663] = 3'b110;
        rom_memory[4664] = 3'b110;
        rom_memory[4665] = 3'b110;
        rom_memory[4666] = 3'b110;
        rom_memory[4667] = 3'b110;
        rom_memory[4668] = 3'b110;
        rom_memory[4669] = 3'b110;
        rom_memory[4670] = 3'b110;
        rom_memory[4671] = 3'b110;
        rom_memory[4672] = 3'b110;
        rom_memory[4673] = 3'b110;
        rom_memory[4674] = 3'b110;
        rom_memory[4675] = 3'b110;
        rom_memory[4676] = 3'b110;
        rom_memory[4677] = 3'b110;
        rom_memory[4678] = 3'b110;
        rom_memory[4679] = 3'b110;
        rom_memory[4680] = 3'b110;
        rom_memory[4681] = 3'b110;
        rom_memory[4682] = 3'b110;
        rom_memory[4683] = 3'b110;
        rom_memory[4684] = 3'b110;
        rom_memory[4685] = 3'b110;
        rom_memory[4686] = 3'b110;
        rom_memory[4687] = 3'b110;
        rom_memory[4688] = 3'b110;
        rom_memory[4689] = 3'b110;
        rom_memory[4690] = 3'b110;
        rom_memory[4691] = 3'b110;
        rom_memory[4692] = 3'b110;
        rom_memory[4693] = 3'b110;
        rom_memory[4694] = 3'b110;
        rom_memory[4695] = 3'b110;
        rom_memory[4696] = 3'b110;
        rom_memory[4697] = 3'b110;
        rom_memory[4698] = 3'b110;
        rom_memory[4699] = 3'b110;
        rom_memory[4700] = 3'b110;
        rom_memory[4701] = 3'b110;
        rom_memory[4702] = 3'b110;
        rom_memory[4703] = 3'b110;
        rom_memory[4704] = 3'b110;
        rom_memory[4705] = 3'b110;
        rom_memory[4706] = 3'b110;
        rom_memory[4707] = 3'b110;
        rom_memory[4708] = 3'b110;
        rom_memory[4709] = 3'b110;
        rom_memory[4710] = 3'b110;
        rom_memory[4711] = 3'b110;
        rom_memory[4712] = 3'b110;
        rom_memory[4713] = 3'b110;
        rom_memory[4714] = 3'b110;
        rom_memory[4715] = 3'b110;
        rom_memory[4716] = 3'b110;
        rom_memory[4717] = 3'b110;
        rom_memory[4718] = 3'b110;
        rom_memory[4719] = 3'b110;
        rom_memory[4720] = 3'b110;
        rom_memory[4721] = 3'b110;
        rom_memory[4722] = 3'b110;
        rom_memory[4723] = 3'b110;
        rom_memory[4724] = 3'b110;
        rom_memory[4725] = 3'b110;
        rom_memory[4726] = 3'b110;
        rom_memory[4727] = 3'b110;
        rom_memory[4728] = 3'b110;
        rom_memory[4729] = 3'b110;
        rom_memory[4730] = 3'b110;
        rom_memory[4731] = 3'b110;
        rom_memory[4732] = 3'b110;
        rom_memory[4733] = 3'b110;
        rom_memory[4734] = 3'b110;
        rom_memory[4735] = 3'b110;
        rom_memory[4736] = 3'b110;
        rom_memory[4737] = 3'b110;
        rom_memory[4738] = 3'b110;
        rom_memory[4739] = 3'b110;
        rom_memory[4740] = 3'b110;
        rom_memory[4741] = 3'b110;
        rom_memory[4742] = 3'b110;
        rom_memory[4743] = 3'b110;
        rom_memory[4744] = 3'b110;
        rom_memory[4745] = 3'b110;
        rom_memory[4746] = 3'b110;
        rom_memory[4747] = 3'b110;
        rom_memory[4748] = 3'b110;
        rom_memory[4749] = 3'b110;
        rom_memory[4750] = 3'b110;
        rom_memory[4751] = 3'b110;
        rom_memory[4752] = 3'b110;
        rom_memory[4753] = 3'b110;
        rom_memory[4754] = 3'b110;
        rom_memory[4755] = 3'b110;
        rom_memory[4756] = 3'b110;
        rom_memory[4757] = 3'b110;
        rom_memory[4758] = 3'b110;
        rom_memory[4759] = 3'b110;
        rom_memory[4760] = 3'b110;
        rom_memory[4761] = 3'b110;
        rom_memory[4762] = 3'b110;
        rom_memory[4763] = 3'b110;
        rom_memory[4764] = 3'b110;
        rom_memory[4765] = 3'b110;
        rom_memory[4766] = 3'b110;
        rom_memory[4767] = 3'b110;
        rom_memory[4768] = 3'b110;
        rom_memory[4769] = 3'b110;
        rom_memory[4770] = 3'b110;
        rom_memory[4771] = 3'b110;
        rom_memory[4772] = 3'b110;
        rom_memory[4773] = 3'b110;
        rom_memory[4774] = 3'b110;
        rom_memory[4775] = 3'b110;
        rom_memory[4776] = 3'b110;
        rom_memory[4777] = 3'b110;
        rom_memory[4778] = 3'b110;
        rom_memory[4779] = 3'b110;
        rom_memory[4780] = 3'b110;
        rom_memory[4781] = 3'b110;
        rom_memory[4782] = 3'b110;
        rom_memory[4783] = 3'b110;
        rom_memory[4784] = 3'b110;
        rom_memory[4785] = 3'b110;
        rom_memory[4786] = 3'b110;
        rom_memory[4787] = 3'b110;
        rom_memory[4788] = 3'b110;
        rom_memory[4789] = 3'b110;
        rom_memory[4790] = 3'b110;
        rom_memory[4791] = 3'b110;
        rom_memory[4792] = 3'b110;
        rom_memory[4793] = 3'b110;
        rom_memory[4794] = 3'b110;
        rom_memory[4795] = 3'b110;
        rom_memory[4796] = 3'b110;
        rom_memory[4797] = 3'b110;
        rom_memory[4798] = 3'b110;
        rom_memory[4799] = 3'b110;
        rom_memory[4800] = 3'b110;
        rom_memory[4801] = 3'b110;
        rom_memory[4802] = 3'b110;
        rom_memory[4803] = 3'b110;
        rom_memory[4804] = 3'b110;
        rom_memory[4805] = 3'b110;
        rom_memory[4806] = 3'b110;
        rom_memory[4807] = 3'b110;
        rom_memory[4808] = 3'b110;
        rom_memory[4809] = 3'b110;
        rom_memory[4810] = 3'b110;
        rom_memory[4811] = 3'b110;
        rom_memory[4812] = 3'b110;
        rom_memory[4813] = 3'b110;
        rom_memory[4814] = 3'b110;
        rom_memory[4815] = 3'b110;
        rom_memory[4816] = 3'b111;
        rom_memory[4817] = 3'b111;
        rom_memory[4818] = 3'b111;
        rom_memory[4819] = 3'b111;
        rom_memory[4820] = 3'b111;
        rom_memory[4821] = 3'b111;
        rom_memory[4822] = 3'b111;
        rom_memory[4823] = 3'b111;
        rom_memory[4824] = 3'b111;
        rom_memory[4825] = 3'b111;
        rom_memory[4826] = 3'b111;
        rom_memory[4827] = 3'b111;
        rom_memory[4828] = 3'b111;
        rom_memory[4829] = 3'b111;
        rom_memory[4830] = 3'b111;
        rom_memory[4831] = 3'b111;
        rom_memory[4832] = 3'b111;
        rom_memory[4833] = 3'b111;
        rom_memory[4834] = 3'b111;
        rom_memory[4835] = 3'b110;
        rom_memory[4836] = 3'b110;
        rom_memory[4837] = 3'b110;
        rom_memory[4838] = 3'b110;
        rom_memory[4839] = 3'b110;
        rom_memory[4840] = 3'b110;
        rom_memory[4841] = 3'b110;
        rom_memory[4842] = 3'b110;
        rom_memory[4843] = 3'b110;
        rom_memory[4844] = 3'b110;
        rom_memory[4845] = 3'b110;
        rom_memory[4846] = 3'b110;
        rom_memory[4847] = 3'b110;
        rom_memory[4848] = 3'b110;
        rom_memory[4849] = 3'b110;
        rom_memory[4850] = 3'b110;
        rom_memory[4851] = 3'b110;
        rom_memory[4852] = 3'b110;
        rom_memory[4853] = 3'b110;
        rom_memory[4854] = 3'b110;
        rom_memory[4855] = 3'b110;
        rom_memory[4856] = 3'b110;
        rom_memory[4857] = 3'b110;
        rom_memory[4858] = 3'b111;
        rom_memory[4859] = 3'b111;
        rom_memory[4860] = 3'b111;
        rom_memory[4861] = 3'b111;
        rom_memory[4862] = 3'b111;
        rom_memory[4863] = 3'b111;
        rom_memory[4864] = 3'b111;
        rom_memory[4865] = 3'b111;
        rom_memory[4866] = 3'b111;
        rom_memory[4867] = 3'b111;
        rom_memory[4868] = 3'b111;
        rom_memory[4869] = 3'b111;
        rom_memory[4870] = 3'b111;
        rom_memory[4871] = 3'b111;
        rom_memory[4872] = 3'b111;
        rom_memory[4873] = 3'b111;
        rom_memory[4874] = 3'b111;
        rom_memory[4875] = 3'b111;
        rom_memory[4876] = 3'b110;
        rom_memory[4877] = 3'b110;
        rom_memory[4878] = 3'b110;
        rom_memory[4879] = 3'b110;
        rom_memory[4880] = 3'b110;
        rom_memory[4881] = 3'b110;
        rom_memory[4882] = 3'b110;
        rom_memory[4883] = 3'b110;
        rom_memory[4884] = 3'b110;
        rom_memory[4885] = 3'b110;
        rom_memory[4886] = 3'b110;
        rom_memory[4887] = 3'b110;
        rom_memory[4888] = 3'b110;
        rom_memory[4889] = 3'b110;
        rom_memory[4890] = 3'b110;
        rom_memory[4891] = 3'b110;
        rom_memory[4892] = 3'b110;
        rom_memory[4893] = 3'b110;
        rom_memory[4894] = 3'b110;
        rom_memory[4895] = 3'b110;
        rom_memory[4896] = 3'b110;
        rom_memory[4897] = 3'b110;
        rom_memory[4898] = 3'b110;
        rom_memory[4899] = 3'b110;
        rom_memory[4900] = 3'b110;
        rom_memory[4901] = 3'b110;
        rom_memory[4902] = 3'b110;
        rom_memory[4903] = 3'b110;
        rom_memory[4904] = 3'b110;
        rom_memory[4905] = 3'b110;
        rom_memory[4906] = 3'b110;
        rom_memory[4907] = 3'b110;
        rom_memory[4908] = 3'b110;
        rom_memory[4909] = 3'b110;
        rom_memory[4910] = 3'b110;
        rom_memory[4911] = 3'b110;
        rom_memory[4912] = 3'b110;
        rom_memory[4913] = 3'b110;
        rom_memory[4914] = 3'b110;
        rom_memory[4915] = 3'b110;
        rom_memory[4916] = 3'b110;
        rom_memory[4917] = 3'b110;
        rom_memory[4918] = 3'b110;
        rom_memory[4919] = 3'b110;
        rom_memory[4920] = 3'b110;
        rom_memory[4921] = 3'b110;
        rom_memory[4922] = 3'b110;
        rom_memory[4923] = 3'b110;
        rom_memory[4924] = 3'b110;
        rom_memory[4925] = 3'b110;
        rom_memory[4926] = 3'b110;
        rom_memory[4927] = 3'b110;
        rom_memory[4928] = 3'b110;
        rom_memory[4929] = 3'b110;
        rom_memory[4930] = 3'b110;
        rom_memory[4931] = 3'b110;
        rom_memory[4932] = 3'b110;
        rom_memory[4933] = 3'b110;
        rom_memory[4934] = 3'b110;
        rom_memory[4935] = 3'b110;
        rom_memory[4936] = 3'b110;
        rom_memory[4937] = 3'b110;
        rom_memory[4938] = 3'b110;
        rom_memory[4939] = 3'b110;
        rom_memory[4940] = 3'b110;
        rom_memory[4941] = 3'b110;
        rom_memory[4942] = 3'b110;
        rom_memory[4943] = 3'b110;
        rom_memory[4944] = 3'b110;
        rom_memory[4945] = 3'b110;
        rom_memory[4946] = 3'b110;
        rom_memory[4947] = 3'b110;
        rom_memory[4948] = 3'b110;
        rom_memory[4949] = 3'b110;
        rom_memory[4950] = 3'b110;
        rom_memory[4951] = 3'b110;
        rom_memory[4952] = 3'b110;
        rom_memory[4953] = 3'b110;
        rom_memory[4954] = 3'b110;
        rom_memory[4955] = 3'b110;
        rom_memory[4956] = 3'b110;
        rom_memory[4957] = 3'b110;
        rom_memory[4958] = 3'b110;
        rom_memory[4959] = 3'b110;
        rom_memory[4960] = 3'b110;
        rom_memory[4961] = 3'b110;
        rom_memory[4962] = 3'b110;
        rom_memory[4963] = 3'b110;
        rom_memory[4964] = 3'b110;
        rom_memory[4965] = 3'b110;
        rom_memory[4966] = 3'b110;
        rom_memory[4967] = 3'b110;
        rom_memory[4968] = 3'b110;
        rom_memory[4969] = 3'b110;
        rom_memory[4970] = 3'b110;
        rom_memory[4971] = 3'b110;
        rom_memory[4972] = 3'b110;
        rom_memory[4973] = 3'b110;
        rom_memory[4974] = 3'b110;
        rom_memory[4975] = 3'b110;
        rom_memory[4976] = 3'b110;
        rom_memory[4977] = 3'b110;
        rom_memory[4978] = 3'b110;
        rom_memory[4979] = 3'b110;
        rom_memory[4980] = 3'b110;
        rom_memory[4981] = 3'b110;
        rom_memory[4982] = 3'b110;
        rom_memory[4983] = 3'b110;
        rom_memory[4984] = 3'b110;
        rom_memory[4985] = 3'b110;
        rom_memory[4986] = 3'b110;
        rom_memory[4987] = 3'b110;
        rom_memory[4988] = 3'b110;
        rom_memory[4989] = 3'b110;
        rom_memory[4990] = 3'b110;
        rom_memory[4991] = 3'b110;
        rom_memory[4992] = 3'b110;
        rom_memory[4993] = 3'b110;
        rom_memory[4994] = 3'b110;
        rom_memory[4995] = 3'b110;
        rom_memory[4996] = 3'b110;
        rom_memory[4997] = 3'b110;
        rom_memory[4998] = 3'b110;
        rom_memory[4999] = 3'b110;
        rom_memory[5000] = 3'b110;
        rom_memory[5001] = 3'b110;
        rom_memory[5002] = 3'b110;
        rom_memory[5003] = 3'b110;
        rom_memory[5004] = 3'b110;
        rom_memory[5005] = 3'b110;
        rom_memory[5006] = 3'b110;
        rom_memory[5007] = 3'b110;
        rom_memory[5008] = 3'b110;
        rom_memory[5009] = 3'b110;
        rom_memory[5010] = 3'b110;
        rom_memory[5011] = 3'b110;
        rom_memory[5012] = 3'b110;
        rom_memory[5013] = 3'b110;
        rom_memory[5014] = 3'b110;
        rom_memory[5015] = 3'b110;
        rom_memory[5016] = 3'b110;
        rom_memory[5017] = 3'b110;
        rom_memory[5018] = 3'b110;
        rom_memory[5019] = 3'b110;
        rom_memory[5020] = 3'b110;
        rom_memory[5021] = 3'b110;
        rom_memory[5022] = 3'b110;
        rom_memory[5023] = 3'b110;
        rom_memory[5024] = 3'b110;
        rom_memory[5025] = 3'b110;
        rom_memory[5026] = 3'b110;
        rom_memory[5027] = 3'b110;
        rom_memory[5028] = 3'b110;
        rom_memory[5029] = 3'b110;
        rom_memory[5030] = 3'b110;
        rom_memory[5031] = 3'b110;
        rom_memory[5032] = 3'b110;
        rom_memory[5033] = 3'b110;
        rom_memory[5034] = 3'b110;
        rom_memory[5035] = 3'b110;
        rom_memory[5036] = 3'b110;
        rom_memory[5037] = 3'b110;
        rom_memory[5038] = 3'b110;
        rom_memory[5039] = 3'b110;
        rom_memory[5040] = 3'b110;
        rom_memory[5041] = 3'b110;
        rom_memory[5042] = 3'b110;
        rom_memory[5043] = 3'b110;
        rom_memory[5044] = 3'b110;
        rom_memory[5045] = 3'b110;
        rom_memory[5046] = 3'b110;
        rom_memory[5047] = 3'b110;
        rom_memory[5048] = 3'b110;
        rom_memory[5049] = 3'b110;
        rom_memory[5050] = 3'b110;
        rom_memory[5051] = 3'b110;
        rom_memory[5052] = 3'b110;
        rom_memory[5053] = 3'b110;
        rom_memory[5054] = 3'b111;
        rom_memory[5055] = 3'b111;
        rom_memory[5056] = 3'b111;
        rom_memory[5057] = 3'b111;
        rom_memory[5058] = 3'b111;
        rom_memory[5059] = 3'b000;
        rom_memory[5060] = 3'b000;
        rom_memory[5061] = 3'b000;
        rom_memory[5062] = 3'b000;
        rom_memory[5063] = 3'b001;
        rom_memory[5064] = 3'b001;
        rom_memory[5065] = 3'b111;
        rom_memory[5066] = 3'b111;
        rom_memory[5067] = 3'b111;
        rom_memory[5068] = 3'b111;
        rom_memory[5069] = 3'b111;
        rom_memory[5070] = 3'b111;
        rom_memory[5071] = 3'b111;
        rom_memory[5072] = 3'b111;
        rom_memory[5073] = 3'b111;
        rom_memory[5074] = 3'b111;
        rom_memory[5075] = 3'b111;
        rom_memory[5076] = 3'b111;
        rom_memory[5077] = 3'b111;
        rom_memory[5078] = 3'b110;
        rom_memory[5079] = 3'b110;
        rom_memory[5080] = 3'b110;
        rom_memory[5081] = 3'b110;
        rom_memory[5082] = 3'b110;
        rom_memory[5083] = 3'b110;
        rom_memory[5084] = 3'b110;
        rom_memory[5085] = 3'b110;
        rom_memory[5086] = 3'b110;
        rom_memory[5087] = 3'b110;
        rom_memory[5088] = 3'b110;
        rom_memory[5089] = 3'b110;
        rom_memory[5090] = 3'b110;
        rom_memory[5091] = 3'b110;
        rom_memory[5092] = 3'b110;
        rom_memory[5093] = 3'b110;
        rom_memory[5094] = 3'b110;
        rom_memory[5095] = 3'b110;
        rom_memory[5096] = 3'b111;
        rom_memory[5097] = 3'b111;
        rom_memory[5098] = 3'b111;
        rom_memory[5099] = 3'b111;
        rom_memory[5100] = 3'b111;
        rom_memory[5101] = 3'b001;
        rom_memory[5102] = 3'b011;
        rom_memory[5103] = 3'b011;
        rom_memory[5104] = 3'b011;
        rom_memory[5105] = 3'b011;
        rom_memory[5106] = 3'b001;
        rom_memory[5107] = 3'b001;
        rom_memory[5108] = 3'b011;
        rom_memory[5109] = 3'b011;
        rom_memory[5110] = 3'b011;
        rom_memory[5111] = 3'b011;
        rom_memory[5112] = 3'b011;
        rom_memory[5113] = 3'b111;
        rom_memory[5114] = 3'b111;
        rom_memory[5115] = 3'b111;
        rom_memory[5116] = 3'b111;
        rom_memory[5117] = 3'b111;
        rom_memory[5118] = 3'b110;
        rom_memory[5119] = 3'b110;
        rom_memory[5120] = 3'b110;
        rom_memory[5121] = 3'b110;
        rom_memory[5122] = 3'b110;
        rom_memory[5123] = 3'b110;
        rom_memory[5124] = 3'b110;
        rom_memory[5125] = 3'b110;
        rom_memory[5126] = 3'b110;
        rom_memory[5127] = 3'b110;
        rom_memory[5128] = 3'b110;
        rom_memory[5129] = 3'b110;
        rom_memory[5130] = 3'b110;
        rom_memory[5131] = 3'b110;
        rom_memory[5132] = 3'b110;
        rom_memory[5133] = 3'b110;
        rom_memory[5134] = 3'b110;
        rom_memory[5135] = 3'b110;
        rom_memory[5136] = 3'b110;
        rom_memory[5137] = 3'b110;
        rom_memory[5138] = 3'b110;
        rom_memory[5139] = 3'b110;
        rom_memory[5140] = 3'b110;
        rom_memory[5141] = 3'b110;
        rom_memory[5142] = 3'b110;
        rom_memory[5143] = 3'b110;
        rom_memory[5144] = 3'b110;
        rom_memory[5145] = 3'b110;
        rom_memory[5146] = 3'b110;
        rom_memory[5147] = 3'b110;
        rom_memory[5148] = 3'b110;
        rom_memory[5149] = 3'b110;
        rom_memory[5150] = 3'b110;
        rom_memory[5151] = 3'b110;
        rom_memory[5152] = 3'b110;
        rom_memory[5153] = 3'b110;
        rom_memory[5154] = 3'b110;
        rom_memory[5155] = 3'b110;
        rom_memory[5156] = 3'b110;
        rom_memory[5157] = 3'b110;
        rom_memory[5158] = 3'b110;
        rom_memory[5159] = 3'b110;
        rom_memory[5160] = 3'b110;
        rom_memory[5161] = 3'b110;
        rom_memory[5162] = 3'b110;
        rom_memory[5163] = 3'b110;
        rom_memory[5164] = 3'b110;
        rom_memory[5165] = 3'b110;
        rom_memory[5166] = 3'b110;
        rom_memory[5167] = 3'b110;
        rom_memory[5168] = 3'b110;
        rom_memory[5169] = 3'b110;
        rom_memory[5170] = 3'b110;
        rom_memory[5171] = 3'b110;
        rom_memory[5172] = 3'b110;
        rom_memory[5173] = 3'b110;
        rom_memory[5174] = 3'b110;
        rom_memory[5175] = 3'b110;
        rom_memory[5176] = 3'b110;
        rom_memory[5177] = 3'b110;
        rom_memory[5178] = 3'b110;
        rom_memory[5179] = 3'b110;
        rom_memory[5180] = 3'b110;
        rom_memory[5181] = 3'b110;
        rom_memory[5182] = 3'b110;
        rom_memory[5183] = 3'b110;
        rom_memory[5184] = 3'b110;
        rom_memory[5185] = 3'b110;
        rom_memory[5186] = 3'b110;
        rom_memory[5187] = 3'b110;
        rom_memory[5188] = 3'b110;
        rom_memory[5189] = 3'b110;
        rom_memory[5190] = 3'b110;
        rom_memory[5191] = 3'b110;
        rom_memory[5192] = 3'b110;
        rom_memory[5193] = 3'b110;
        rom_memory[5194] = 3'b110;
        rom_memory[5195] = 3'b110;
        rom_memory[5196] = 3'b110;
        rom_memory[5197] = 3'b110;
        rom_memory[5198] = 3'b110;
        rom_memory[5199] = 3'b110;
        rom_memory[5200] = 3'b110;
        rom_memory[5201] = 3'b110;
        rom_memory[5202] = 3'b110;
        rom_memory[5203] = 3'b110;
        rom_memory[5204] = 3'b110;
        rom_memory[5205] = 3'b110;
        rom_memory[5206] = 3'b110;
        rom_memory[5207] = 3'b110;
        rom_memory[5208] = 3'b110;
        rom_memory[5209] = 3'b110;
        rom_memory[5210] = 3'b110;
        rom_memory[5211] = 3'b110;
        rom_memory[5212] = 3'b110;
        rom_memory[5213] = 3'b110;
        rom_memory[5214] = 3'b110;
        rom_memory[5215] = 3'b110;
        rom_memory[5216] = 3'b110;
        rom_memory[5217] = 3'b110;
        rom_memory[5218] = 3'b110;
        rom_memory[5219] = 3'b110;
        rom_memory[5220] = 3'b110;
        rom_memory[5221] = 3'b110;
        rom_memory[5222] = 3'b110;
        rom_memory[5223] = 3'b110;
        rom_memory[5224] = 3'b110;
        rom_memory[5225] = 3'b110;
        rom_memory[5226] = 3'b110;
        rom_memory[5227] = 3'b110;
        rom_memory[5228] = 3'b110;
        rom_memory[5229] = 3'b110;
        rom_memory[5230] = 3'b110;
        rom_memory[5231] = 3'b110;
        rom_memory[5232] = 3'b110;
        rom_memory[5233] = 3'b110;
        rom_memory[5234] = 3'b110;
        rom_memory[5235] = 3'b110;
        rom_memory[5236] = 3'b110;
        rom_memory[5237] = 3'b110;
        rom_memory[5238] = 3'b110;
        rom_memory[5239] = 3'b110;
        rom_memory[5240] = 3'b110;
        rom_memory[5241] = 3'b110;
        rom_memory[5242] = 3'b110;
        rom_memory[5243] = 3'b110;
        rom_memory[5244] = 3'b110;
        rom_memory[5245] = 3'b110;
        rom_memory[5246] = 3'b110;
        rom_memory[5247] = 3'b110;
        rom_memory[5248] = 3'b110;
        rom_memory[5249] = 3'b110;
        rom_memory[5250] = 3'b110;
        rom_memory[5251] = 3'b110;
        rom_memory[5252] = 3'b110;
        rom_memory[5253] = 3'b110;
        rom_memory[5254] = 3'b110;
        rom_memory[5255] = 3'b110;
        rom_memory[5256] = 3'b110;
        rom_memory[5257] = 3'b110;
        rom_memory[5258] = 3'b110;
        rom_memory[5259] = 3'b110;
        rom_memory[5260] = 3'b110;
        rom_memory[5261] = 3'b110;
        rom_memory[5262] = 3'b110;
        rom_memory[5263] = 3'b110;
        rom_memory[5264] = 3'b110;
        rom_memory[5265] = 3'b110;
        rom_memory[5266] = 3'b110;
        rom_memory[5267] = 3'b110;
        rom_memory[5268] = 3'b110;
        rom_memory[5269] = 3'b110;
        rom_memory[5270] = 3'b110;
        rom_memory[5271] = 3'b110;
        rom_memory[5272] = 3'b110;
        rom_memory[5273] = 3'b110;
        rom_memory[5274] = 3'b110;
        rom_memory[5275] = 3'b110;
        rom_memory[5276] = 3'b110;
        rom_memory[5277] = 3'b110;
        rom_memory[5278] = 3'b110;
        rom_memory[5279] = 3'b110;
        rom_memory[5280] = 3'b110;
        rom_memory[5281] = 3'b110;
        rom_memory[5282] = 3'b110;
        rom_memory[5283] = 3'b110;
        rom_memory[5284] = 3'b110;
        rom_memory[5285] = 3'b110;
        rom_memory[5286] = 3'b110;
        rom_memory[5287] = 3'b110;
        rom_memory[5288] = 3'b110;
        rom_memory[5289] = 3'b110;
        rom_memory[5290] = 3'b110;
        rom_memory[5291] = 3'b110;
        rom_memory[5292] = 3'b111;
        rom_memory[5293] = 3'b111;
        rom_memory[5294] = 3'b111;
        rom_memory[5295] = 3'b111;
        rom_memory[5296] = 3'b100;
        rom_memory[5297] = 3'b100;
        rom_memory[5298] = 3'b000;
        rom_memory[5299] = 3'b000;
        rom_memory[5300] = 3'b000;
        rom_memory[5301] = 3'b000;
        rom_memory[5302] = 3'b000;
        rom_memory[5303] = 3'b000;
        rom_memory[5304] = 3'b000;
        rom_memory[5305] = 3'b000;
        rom_memory[5306] = 3'b000;
        rom_memory[5307] = 3'b000;
        rom_memory[5308] = 3'b000;
        rom_memory[5309] = 3'b000;
        rom_memory[5310] = 3'b000;
        rom_memory[5311] = 3'b000;
        rom_memory[5312] = 3'b111;
        rom_memory[5313] = 3'b111;
        rom_memory[5314] = 3'b111;
        rom_memory[5315] = 3'b111;
        rom_memory[5316] = 3'b111;
        rom_memory[5317] = 3'b111;
        rom_memory[5318] = 3'b111;
        rom_memory[5319] = 3'b111;
        rom_memory[5320] = 3'b110;
        rom_memory[5321] = 3'b110;
        rom_memory[5322] = 3'b110;
        rom_memory[5323] = 3'b110;
        rom_memory[5324] = 3'b110;
        rom_memory[5325] = 3'b110;
        rom_memory[5326] = 3'b110;
        rom_memory[5327] = 3'b110;
        rom_memory[5328] = 3'b110;
        rom_memory[5329] = 3'b110;
        rom_memory[5330] = 3'b110;
        rom_memory[5331] = 3'b110;
        rom_memory[5332] = 3'b110;
        rom_memory[5333] = 3'b110;
        rom_memory[5334] = 3'b110;
        rom_memory[5335] = 3'b111;
        rom_memory[5336] = 3'b111;
        rom_memory[5337] = 3'b001;
        rom_memory[5338] = 3'b011;
        rom_memory[5339] = 3'b011;
        rom_memory[5340] = 3'b001;
        rom_memory[5341] = 3'b001;
        rom_memory[5342] = 3'b011;
        rom_memory[5343] = 3'b001;
        rom_memory[5344] = 3'b001;
        rom_memory[5345] = 3'b001;
        rom_memory[5346] = 3'b000;
        rom_memory[5347] = 3'b001;
        rom_memory[5348] = 3'b011;
        rom_memory[5349] = 3'b001;
        rom_memory[5350] = 3'b011;
        rom_memory[5351] = 3'b011;
        rom_memory[5352] = 3'b011;
        rom_memory[5353] = 3'b011;
        rom_memory[5354] = 3'b111;
        rom_memory[5355] = 3'b111;
        rom_memory[5356] = 3'b111;
        rom_memory[5357] = 3'b111;
        rom_memory[5358] = 3'b111;
        rom_memory[5359] = 3'b111;
        rom_memory[5360] = 3'b110;
        rom_memory[5361] = 3'b110;
        rom_memory[5362] = 3'b110;
        rom_memory[5363] = 3'b110;
        rom_memory[5364] = 3'b110;
        rom_memory[5365] = 3'b110;
        rom_memory[5366] = 3'b110;
        rom_memory[5367] = 3'b110;
        rom_memory[5368] = 3'b110;
        rom_memory[5369] = 3'b110;
        rom_memory[5370] = 3'b110;
        rom_memory[5371] = 3'b110;
        rom_memory[5372] = 3'b110;
        rom_memory[5373] = 3'b110;
        rom_memory[5374] = 3'b110;
        rom_memory[5375] = 3'b110;
        rom_memory[5376] = 3'b110;
        rom_memory[5377] = 3'b110;
        rom_memory[5378] = 3'b110;
        rom_memory[5379] = 3'b110;
        rom_memory[5380] = 3'b110;
        rom_memory[5381] = 3'b110;
        rom_memory[5382] = 3'b110;
        rom_memory[5383] = 3'b110;
        rom_memory[5384] = 3'b110;
        rom_memory[5385] = 3'b110;
        rom_memory[5386] = 3'b110;
        rom_memory[5387] = 3'b110;
        rom_memory[5388] = 3'b110;
        rom_memory[5389] = 3'b110;
        rom_memory[5390] = 3'b110;
        rom_memory[5391] = 3'b110;
        rom_memory[5392] = 3'b110;
        rom_memory[5393] = 3'b110;
        rom_memory[5394] = 3'b110;
        rom_memory[5395] = 3'b110;
        rom_memory[5396] = 3'b110;
        rom_memory[5397] = 3'b110;
        rom_memory[5398] = 3'b110;
        rom_memory[5399] = 3'b110;
        rom_memory[5400] = 3'b110;
        rom_memory[5401] = 3'b110;
        rom_memory[5402] = 3'b110;
        rom_memory[5403] = 3'b110;
        rom_memory[5404] = 3'b110;
        rom_memory[5405] = 3'b110;
        rom_memory[5406] = 3'b110;
        rom_memory[5407] = 3'b110;
        rom_memory[5408] = 3'b110;
        rom_memory[5409] = 3'b110;
        rom_memory[5410] = 3'b110;
        rom_memory[5411] = 3'b110;
        rom_memory[5412] = 3'b110;
        rom_memory[5413] = 3'b110;
        rom_memory[5414] = 3'b110;
        rom_memory[5415] = 3'b110;
        rom_memory[5416] = 3'b110;
        rom_memory[5417] = 3'b110;
        rom_memory[5418] = 3'b110;
        rom_memory[5419] = 3'b110;
        rom_memory[5420] = 3'b110;
        rom_memory[5421] = 3'b110;
        rom_memory[5422] = 3'b110;
        rom_memory[5423] = 3'b110;
        rom_memory[5424] = 3'b110;
        rom_memory[5425] = 3'b110;
        rom_memory[5426] = 3'b110;
        rom_memory[5427] = 3'b110;
        rom_memory[5428] = 3'b110;
        rom_memory[5429] = 3'b110;
        rom_memory[5430] = 3'b110;
        rom_memory[5431] = 3'b110;
        rom_memory[5432] = 3'b110;
        rom_memory[5433] = 3'b110;
        rom_memory[5434] = 3'b110;
        rom_memory[5435] = 3'b110;
        rom_memory[5436] = 3'b110;
        rom_memory[5437] = 3'b110;
        rom_memory[5438] = 3'b110;
        rom_memory[5439] = 3'b110;
        rom_memory[5440] = 3'b110;
        rom_memory[5441] = 3'b110;
        rom_memory[5442] = 3'b110;
        rom_memory[5443] = 3'b110;
        rom_memory[5444] = 3'b110;
        rom_memory[5445] = 3'b110;
        rom_memory[5446] = 3'b110;
        rom_memory[5447] = 3'b110;
        rom_memory[5448] = 3'b110;
        rom_memory[5449] = 3'b110;
        rom_memory[5450] = 3'b110;
        rom_memory[5451] = 3'b110;
        rom_memory[5452] = 3'b110;
        rom_memory[5453] = 3'b110;
        rom_memory[5454] = 3'b110;
        rom_memory[5455] = 3'b110;
        rom_memory[5456] = 3'b110;
        rom_memory[5457] = 3'b110;
        rom_memory[5458] = 3'b110;
        rom_memory[5459] = 3'b110;
        rom_memory[5460] = 3'b110;
        rom_memory[5461] = 3'b110;
        rom_memory[5462] = 3'b110;
        rom_memory[5463] = 3'b110;
        rom_memory[5464] = 3'b110;
        rom_memory[5465] = 3'b110;
        rom_memory[5466] = 3'b110;
        rom_memory[5467] = 3'b110;
        rom_memory[5468] = 3'b110;
        rom_memory[5469] = 3'b110;
        rom_memory[5470] = 3'b110;
        rom_memory[5471] = 3'b110;
        rom_memory[5472] = 3'b110;
        rom_memory[5473] = 3'b110;
        rom_memory[5474] = 3'b110;
        rom_memory[5475] = 3'b110;
        rom_memory[5476] = 3'b110;
        rom_memory[5477] = 3'b110;
        rom_memory[5478] = 3'b110;
        rom_memory[5479] = 3'b110;
        rom_memory[5480] = 3'b110;
        rom_memory[5481] = 3'b110;
        rom_memory[5482] = 3'b110;
        rom_memory[5483] = 3'b110;
        rom_memory[5484] = 3'b110;
        rom_memory[5485] = 3'b110;
        rom_memory[5486] = 3'b110;
        rom_memory[5487] = 3'b110;
        rom_memory[5488] = 3'b110;
        rom_memory[5489] = 3'b110;
        rom_memory[5490] = 3'b110;
        rom_memory[5491] = 3'b110;
        rom_memory[5492] = 3'b110;
        rom_memory[5493] = 3'b110;
        rom_memory[5494] = 3'b110;
        rom_memory[5495] = 3'b110;
        rom_memory[5496] = 3'b110;
        rom_memory[5497] = 3'b110;
        rom_memory[5498] = 3'b110;
        rom_memory[5499] = 3'b110;
        rom_memory[5500] = 3'b110;
        rom_memory[5501] = 3'b110;
        rom_memory[5502] = 3'b110;
        rom_memory[5503] = 3'b110;
        rom_memory[5504] = 3'b110;
        rom_memory[5505] = 3'b110;
        rom_memory[5506] = 3'b110;
        rom_memory[5507] = 3'b110;
        rom_memory[5508] = 3'b110;
        rom_memory[5509] = 3'b110;
        rom_memory[5510] = 3'b110;
        rom_memory[5511] = 3'b110;
        rom_memory[5512] = 3'b110;
        rom_memory[5513] = 3'b110;
        rom_memory[5514] = 3'b110;
        rom_memory[5515] = 3'b110;
        rom_memory[5516] = 3'b110;
        rom_memory[5517] = 3'b110;
        rom_memory[5518] = 3'b110;
        rom_memory[5519] = 3'b110;
        rom_memory[5520] = 3'b110;
        rom_memory[5521] = 3'b110;
        rom_memory[5522] = 3'b110;
        rom_memory[5523] = 3'b110;
        rom_memory[5524] = 3'b110;
        rom_memory[5525] = 3'b110;
        rom_memory[5526] = 3'b110;
        rom_memory[5527] = 3'b110;
        rom_memory[5528] = 3'b110;
        rom_memory[5529] = 3'b110;
        rom_memory[5530] = 3'b110;
        rom_memory[5531] = 3'b111;
        rom_memory[5532] = 3'b111;
        rom_memory[5533] = 3'b111;
        rom_memory[5534] = 3'b110;
        rom_memory[5535] = 3'b110;
        rom_memory[5536] = 3'b110;
        rom_memory[5537] = 3'b110;
        rom_memory[5538] = 3'b110;
        rom_memory[5539] = 3'b110;
        rom_memory[5540] = 3'b110;
        rom_memory[5541] = 3'b110;
        rom_memory[5542] = 3'b110;
        rom_memory[5543] = 3'b100;
        rom_memory[5544] = 3'b000;
        rom_memory[5545] = 3'b000;
        rom_memory[5546] = 3'b000;
        rom_memory[5547] = 3'b000;
        rom_memory[5548] = 3'b000;
        rom_memory[5549] = 3'b000;
        rom_memory[5550] = 3'b000;
        rom_memory[5551] = 3'b000;
        rom_memory[5552] = 3'b000;
        rom_memory[5553] = 3'b000;
        rom_memory[5554] = 3'b000;
        rom_memory[5555] = 3'b111;
        rom_memory[5556] = 3'b111;
        rom_memory[5557] = 3'b111;
        rom_memory[5558] = 3'b111;
        rom_memory[5559] = 3'b111;
        rom_memory[5560] = 3'b111;
        rom_memory[5561] = 3'b111;
        rom_memory[5562] = 3'b111;
        rom_memory[5563] = 3'b110;
        rom_memory[5564] = 3'b110;
        rom_memory[5565] = 3'b110;
        rom_memory[5566] = 3'b110;
        rom_memory[5567] = 3'b110;
        rom_memory[5568] = 3'b110;
        rom_memory[5569] = 3'b110;
        rom_memory[5570] = 3'b110;
        rom_memory[5571] = 3'b110;
        rom_memory[5572] = 3'b110;
        rom_memory[5573] = 3'b111;
        rom_memory[5574] = 3'b111;
        rom_memory[5575] = 3'b111;
        rom_memory[5576] = 3'b000;
        rom_memory[5577] = 3'b001;
        rom_memory[5578] = 3'b001;
        rom_memory[5579] = 3'b001;
        rom_memory[5580] = 3'b001;
        rom_memory[5581] = 3'b001;
        rom_memory[5582] = 3'b001;
        rom_memory[5583] = 3'b000;
        rom_memory[5584] = 3'b000;
        rom_memory[5585] = 3'b000;
        rom_memory[5586] = 3'b000;
        rom_memory[5587] = 3'b001;
        rom_memory[5588] = 3'b011;
        rom_memory[5589] = 3'b000;
        rom_memory[5590] = 3'b011;
        rom_memory[5591] = 3'b011;
        rom_memory[5592] = 3'b011;
        rom_memory[5593] = 3'b011;
        rom_memory[5594] = 3'b011;
        rom_memory[5595] = 3'b011;
        rom_memory[5596] = 3'b011;
        rom_memory[5597] = 3'b011;
        rom_memory[5598] = 3'b011;
        rom_memory[5599] = 3'b111;
        rom_memory[5600] = 3'b111;
        rom_memory[5601] = 3'b111;
        rom_memory[5602] = 3'b110;
        rom_memory[5603] = 3'b110;
        rom_memory[5604] = 3'b110;
        rom_memory[5605] = 3'b110;
        rom_memory[5606] = 3'b110;
        rom_memory[5607] = 3'b110;
        rom_memory[5608] = 3'b110;
        rom_memory[5609] = 3'b110;
        rom_memory[5610] = 3'b110;
        rom_memory[5611] = 3'b110;
        rom_memory[5612] = 3'b110;
        rom_memory[5613] = 3'b110;
        rom_memory[5614] = 3'b110;
        rom_memory[5615] = 3'b110;
        rom_memory[5616] = 3'b110;
        rom_memory[5617] = 3'b110;
        rom_memory[5618] = 3'b110;
        rom_memory[5619] = 3'b110;
        rom_memory[5620] = 3'b110;
        rom_memory[5621] = 3'b110;
        rom_memory[5622] = 3'b110;
        rom_memory[5623] = 3'b110;
        rom_memory[5624] = 3'b110;
        rom_memory[5625] = 3'b110;
        rom_memory[5626] = 3'b110;
        rom_memory[5627] = 3'b110;
        rom_memory[5628] = 3'b110;
        rom_memory[5629] = 3'b110;
        rom_memory[5630] = 3'b110;
        rom_memory[5631] = 3'b110;
        rom_memory[5632] = 3'b110;
        rom_memory[5633] = 3'b110;
        rom_memory[5634] = 3'b110;
        rom_memory[5635] = 3'b110;
        rom_memory[5636] = 3'b110;
        rom_memory[5637] = 3'b110;
        rom_memory[5638] = 3'b110;
        rom_memory[5639] = 3'b110;
        rom_memory[5640] = 3'b110;
        rom_memory[5641] = 3'b110;
        rom_memory[5642] = 3'b110;
        rom_memory[5643] = 3'b110;
        rom_memory[5644] = 3'b110;
        rom_memory[5645] = 3'b110;
        rom_memory[5646] = 3'b110;
        rom_memory[5647] = 3'b110;
        rom_memory[5648] = 3'b110;
        rom_memory[5649] = 3'b110;
        rom_memory[5650] = 3'b110;
        rom_memory[5651] = 3'b110;
        rom_memory[5652] = 3'b110;
        rom_memory[5653] = 3'b110;
        rom_memory[5654] = 3'b110;
        rom_memory[5655] = 3'b110;
        rom_memory[5656] = 3'b110;
        rom_memory[5657] = 3'b110;
        rom_memory[5658] = 3'b110;
        rom_memory[5659] = 3'b110;
        rom_memory[5660] = 3'b110;
        rom_memory[5661] = 3'b110;
        rom_memory[5662] = 3'b110;
        rom_memory[5663] = 3'b110;
        rom_memory[5664] = 3'b110;
        rom_memory[5665] = 3'b110;
        rom_memory[5666] = 3'b110;
        rom_memory[5667] = 3'b110;
        rom_memory[5668] = 3'b110;
        rom_memory[5669] = 3'b110;
        rom_memory[5670] = 3'b110;
        rom_memory[5671] = 3'b110;
        rom_memory[5672] = 3'b110;
        rom_memory[5673] = 3'b110;
        rom_memory[5674] = 3'b110;
        rom_memory[5675] = 3'b110;
        rom_memory[5676] = 3'b110;
        rom_memory[5677] = 3'b110;
        rom_memory[5678] = 3'b110;
        rom_memory[5679] = 3'b110;
        rom_memory[5680] = 3'b110;
        rom_memory[5681] = 3'b110;
        rom_memory[5682] = 3'b110;
        rom_memory[5683] = 3'b110;
        rom_memory[5684] = 3'b110;
        rom_memory[5685] = 3'b110;
        rom_memory[5686] = 3'b110;
        rom_memory[5687] = 3'b110;
        rom_memory[5688] = 3'b110;
        rom_memory[5689] = 3'b110;
        rom_memory[5690] = 3'b110;
        rom_memory[5691] = 3'b110;
        rom_memory[5692] = 3'b110;
        rom_memory[5693] = 3'b110;
        rom_memory[5694] = 3'b110;
        rom_memory[5695] = 3'b110;
        rom_memory[5696] = 3'b110;
        rom_memory[5697] = 3'b110;
        rom_memory[5698] = 3'b110;
        rom_memory[5699] = 3'b110;
        rom_memory[5700] = 3'b110;
        rom_memory[5701] = 3'b110;
        rom_memory[5702] = 3'b110;
        rom_memory[5703] = 3'b110;
        rom_memory[5704] = 3'b110;
        rom_memory[5705] = 3'b110;
        rom_memory[5706] = 3'b110;
        rom_memory[5707] = 3'b110;
        rom_memory[5708] = 3'b110;
        rom_memory[5709] = 3'b110;
        rom_memory[5710] = 3'b110;
        rom_memory[5711] = 3'b110;
        rom_memory[5712] = 3'b110;
        rom_memory[5713] = 3'b110;
        rom_memory[5714] = 3'b110;
        rom_memory[5715] = 3'b110;
        rom_memory[5716] = 3'b110;
        rom_memory[5717] = 3'b110;
        rom_memory[5718] = 3'b110;
        rom_memory[5719] = 3'b110;
        rom_memory[5720] = 3'b110;
        rom_memory[5721] = 3'b110;
        rom_memory[5722] = 3'b110;
        rom_memory[5723] = 3'b110;
        rom_memory[5724] = 3'b110;
        rom_memory[5725] = 3'b110;
        rom_memory[5726] = 3'b110;
        rom_memory[5727] = 3'b110;
        rom_memory[5728] = 3'b110;
        rom_memory[5729] = 3'b110;
        rom_memory[5730] = 3'b110;
        rom_memory[5731] = 3'b110;
        rom_memory[5732] = 3'b110;
        rom_memory[5733] = 3'b110;
        rom_memory[5734] = 3'b110;
        rom_memory[5735] = 3'b110;
        rom_memory[5736] = 3'b110;
        rom_memory[5737] = 3'b110;
        rom_memory[5738] = 3'b110;
        rom_memory[5739] = 3'b110;
        rom_memory[5740] = 3'b110;
        rom_memory[5741] = 3'b110;
        rom_memory[5742] = 3'b110;
        rom_memory[5743] = 3'b110;
        rom_memory[5744] = 3'b110;
        rom_memory[5745] = 3'b110;
        rom_memory[5746] = 3'b110;
        rom_memory[5747] = 3'b110;
        rom_memory[5748] = 3'b110;
        rom_memory[5749] = 3'b110;
        rom_memory[5750] = 3'b110;
        rom_memory[5751] = 3'b110;
        rom_memory[5752] = 3'b110;
        rom_memory[5753] = 3'b110;
        rom_memory[5754] = 3'b110;
        rom_memory[5755] = 3'b110;
        rom_memory[5756] = 3'b110;
        rom_memory[5757] = 3'b110;
        rom_memory[5758] = 3'b110;
        rom_memory[5759] = 3'b110;
        rom_memory[5760] = 3'b110;
        rom_memory[5761] = 3'b110;
        rom_memory[5762] = 3'b110;
        rom_memory[5763] = 3'b110;
        rom_memory[5764] = 3'b110;
        rom_memory[5765] = 3'b110;
        rom_memory[5766] = 3'b110;
        rom_memory[5767] = 3'b110;
        rom_memory[5768] = 3'b110;
        rom_memory[5769] = 3'b110;
        rom_memory[5770] = 3'b110;
        rom_memory[5771] = 3'b110;
        rom_memory[5772] = 3'b110;
        rom_memory[5773] = 3'b110;
        rom_memory[5774] = 3'b110;
        rom_memory[5775] = 3'b110;
        rom_memory[5776] = 3'b110;
        rom_memory[5777] = 3'b110;
        rom_memory[5778] = 3'b110;
        rom_memory[5779] = 3'b110;
        rom_memory[5780] = 3'b110;
        rom_memory[5781] = 3'b110;
        rom_memory[5782] = 3'b110;
        rom_memory[5783] = 3'b110;
        rom_memory[5784] = 3'b110;
        rom_memory[5785] = 3'b110;
        rom_memory[5786] = 3'b110;
        rom_memory[5787] = 3'b110;
        rom_memory[5788] = 3'b110;
        rom_memory[5789] = 3'b000;
        rom_memory[5790] = 3'b000;
        rom_memory[5791] = 3'b000;
        rom_memory[5792] = 3'b000;
        rom_memory[5793] = 3'b000;
        rom_memory[5794] = 3'b000;
        rom_memory[5795] = 3'b000;
        rom_memory[5796] = 3'b000;
        rom_memory[5797] = 3'b001;
        rom_memory[5798] = 3'b111;
        rom_memory[5799] = 3'b111;
        rom_memory[5800] = 3'b111;
        rom_memory[5801] = 3'b111;
        rom_memory[5802] = 3'b111;
        rom_memory[5803] = 3'b111;
        rom_memory[5804] = 3'b111;
        rom_memory[5805] = 3'b110;
        rom_memory[5806] = 3'b110;
        rom_memory[5807] = 3'b110;
        rom_memory[5808] = 3'b110;
        rom_memory[5809] = 3'b110;
        rom_memory[5810] = 3'b110;
        rom_memory[5811] = 3'b110;
        rom_memory[5812] = 3'b111;
        rom_memory[5813] = 3'b111;
        rom_memory[5814] = 3'b111;
        rom_memory[5815] = 3'b000;
        rom_memory[5816] = 3'b000;
        rom_memory[5817] = 3'b000;
        rom_memory[5818] = 3'b000;
        rom_memory[5819] = 3'b000;
        rom_memory[5820] = 3'b000;
        rom_memory[5821] = 3'b000;
        rom_memory[5822] = 3'b000;
        rom_memory[5823] = 3'b000;
        rom_memory[5824] = 3'b000;
        rom_memory[5825] = 3'b000;
        rom_memory[5826] = 3'b000;
        rom_memory[5827] = 3'b000;
        rom_memory[5828] = 3'b001;
        rom_memory[5829] = 3'b000;
        rom_memory[5830] = 3'b011;
        rom_memory[5831] = 3'b000;
        rom_memory[5832] = 3'b000;
        rom_memory[5833] = 3'b011;
        rom_memory[5834] = 3'b011;
        rom_memory[5835] = 3'b011;
        rom_memory[5836] = 3'b001;
        rom_memory[5837] = 3'b011;
        rom_memory[5838] = 3'b011;
        rom_memory[5839] = 3'b011;
        rom_memory[5840] = 3'b011;
        rom_memory[5841] = 3'b111;
        rom_memory[5842] = 3'b111;
        rom_memory[5843] = 3'b110;
        rom_memory[5844] = 3'b110;
        rom_memory[5845] = 3'b110;
        rom_memory[5846] = 3'b110;
        rom_memory[5847] = 3'b110;
        rom_memory[5848] = 3'b110;
        rom_memory[5849] = 3'b110;
        rom_memory[5850] = 3'b110;
        rom_memory[5851] = 3'b110;
        rom_memory[5852] = 3'b110;
        rom_memory[5853] = 3'b110;
        rom_memory[5854] = 3'b110;
        rom_memory[5855] = 3'b110;
        rom_memory[5856] = 3'b110;
        rom_memory[5857] = 3'b110;
        rom_memory[5858] = 3'b110;
        rom_memory[5859] = 3'b110;
        rom_memory[5860] = 3'b110;
        rom_memory[5861] = 3'b110;
        rom_memory[5862] = 3'b110;
        rom_memory[5863] = 3'b110;
        rom_memory[5864] = 3'b110;
        rom_memory[5865] = 3'b110;
        rom_memory[5866] = 3'b110;
        rom_memory[5867] = 3'b110;
        rom_memory[5868] = 3'b110;
        rom_memory[5869] = 3'b110;
        rom_memory[5870] = 3'b110;
        rom_memory[5871] = 3'b110;
        rom_memory[5872] = 3'b110;
        rom_memory[5873] = 3'b110;
        rom_memory[5874] = 3'b110;
        rom_memory[5875] = 3'b110;
        rom_memory[5876] = 3'b110;
        rom_memory[5877] = 3'b110;
        rom_memory[5878] = 3'b110;
        rom_memory[5879] = 3'b110;
        rom_memory[5880] = 3'b110;
        rom_memory[5881] = 3'b110;
        rom_memory[5882] = 3'b110;
        rom_memory[5883] = 3'b110;
        rom_memory[5884] = 3'b110;
        rom_memory[5885] = 3'b110;
        rom_memory[5886] = 3'b110;
        rom_memory[5887] = 3'b110;
        rom_memory[5888] = 3'b110;
        rom_memory[5889] = 3'b110;
        rom_memory[5890] = 3'b110;
        rom_memory[5891] = 3'b110;
        rom_memory[5892] = 3'b110;
        rom_memory[5893] = 3'b110;
        rom_memory[5894] = 3'b110;
        rom_memory[5895] = 3'b110;
        rom_memory[5896] = 3'b110;
        rom_memory[5897] = 3'b110;
        rom_memory[5898] = 3'b110;
        rom_memory[5899] = 3'b110;
        rom_memory[5900] = 3'b110;
        rom_memory[5901] = 3'b110;
        rom_memory[5902] = 3'b110;
        rom_memory[5903] = 3'b110;
        rom_memory[5904] = 3'b110;
        rom_memory[5905] = 3'b110;
        rom_memory[5906] = 3'b110;
        rom_memory[5907] = 3'b110;
        rom_memory[5908] = 3'b110;
        rom_memory[5909] = 3'b110;
        rom_memory[5910] = 3'b110;
        rom_memory[5911] = 3'b110;
        rom_memory[5912] = 3'b110;
        rom_memory[5913] = 3'b110;
        rom_memory[5914] = 3'b110;
        rom_memory[5915] = 3'b110;
        rom_memory[5916] = 3'b110;
        rom_memory[5917] = 3'b110;
        rom_memory[5918] = 3'b110;
        rom_memory[5919] = 3'b110;
        rom_memory[5920] = 3'b110;
        rom_memory[5921] = 3'b110;
        rom_memory[5922] = 3'b110;
        rom_memory[5923] = 3'b110;
        rom_memory[5924] = 3'b110;
        rom_memory[5925] = 3'b110;
        rom_memory[5926] = 3'b110;
        rom_memory[5927] = 3'b110;
        rom_memory[5928] = 3'b110;
        rom_memory[5929] = 3'b110;
        rom_memory[5930] = 3'b110;
        rom_memory[5931] = 3'b110;
        rom_memory[5932] = 3'b110;
        rom_memory[5933] = 3'b110;
        rom_memory[5934] = 3'b110;
        rom_memory[5935] = 3'b110;
        rom_memory[5936] = 3'b110;
        rom_memory[5937] = 3'b110;
        rom_memory[5938] = 3'b110;
        rom_memory[5939] = 3'b110;
        rom_memory[5940] = 3'b110;
        rom_memory[5941] = 3'b110;
        rom_memory[5942] = 3'b110;
        rom_memory[5943] = 3'b110;
        rom_memory[5944] = 3'b110;
        rom_memory[5945] = 3'b110;
        rom_memory[5946] = 3'b110;
        rom_memory[5947] = 3'b110;
        rom_memory[5948] = 3'b110;
        rom_memory[5949] = 3'b110;
        rom_memory[5950] = 3'b110;
        rom_memory[5951] = 3'b110;
        rom_memory[5952] = 3'b110;
        rom_memory[5953] = 3'b110;
        rom_memory[5954] = 3'b110;
        rom_memory[5955] = 3'b110;
        rom_memory[5956] = 3'b110;
        rom_memory[5957] = 3'b110;
        rom_memory[5958] = 3'b110;
        rom_memory[5959] = 3'b110;
        rom_memory[5960] = 3'b110;
        rom_memory[5961] = 3'b110;
        rom_memory[5962] = 3'b110;
        rom_memory[5963] = 3'b110;
        rom_memory[5964] = 3'b110;
        rom_memory[5965] = 3'b110;
        rom_memory[5966] = 3'b110;
        rom_memory[5967] = 3'b110;
        rom_memory[5968] = 3'b110;
        rom_memory[5969] = 3'b110;
        rom_memory[5970] = 3'b110;
        rom_memory[5971] = 3'b110;
        rom_memory[5972] = 3'b110;
        rom_memory[5973] = 3'b110;
        rom_memory[5974] = 3'b110;
        rom_memory[5975] = 3'b110;
        rom_memory[5976] = 3'b110;
        rom_memory[5977] = 3'b110;
        rom_memory[5978] = 3'b110;
        rom_memory[5979] = 3'b110;
        rom_memory[5980] = 3'b110;
        rom_memory[5981] = 3'b110;
        rom_memory[5982] = 3'b110;
        rom_memory[5983] = 3'b110;
        rom_memory[5984] = 3'b110;
        rom_memory[5985] = 3'b110;
        rom_memory[5986] = 3'b110;
        rom_memory[5987] = 3'b110;
        rom_memory[5988] = 3'b110;
        rom_memory[5989] = 3'b110;
        rom_memory[5990] = 3'b110;
        rom_memory[5991] = 3'b110;
        rom_memory[5992] = 3'b110;
        rom_memory[5993] = 3'b110;
        rom_memory[5994] = 3'b110;
        rom_memory[5995] = 3'b110;
        rom_memory[5996] = 3'b110;
        rom_memory[5997] = 3'b110;
        rom_memory[5998] = 3'b110;
        rom_memory[5999] = 3'b110;
        rom_memory[6000] = 3'b110;
        rom_memory[6001] = 3'b110;
        rom_memory[6002] = 3'b110;
        rom_memory[6003] = 3'b110;
        rom_memory[6004] = 3'b110;
        rom_memory[6005] = 3'b110;
        rom_memory[6006] = 3'b110;
        rom_memory[6007] = 3'b110;
        rom_memory[6008] = 3'b110;
        rom_memory[6009] = 3'b110;
        rom_memory[6010] = 3'b110;
        rom_memory[6011] = 3'b110;
        rom_memory[6012] = 3'b110;
        rom_memory[6013] = 3'b110;
        rom_memory[6014] = 3'b110;
        rom_memory[6015] = 3'b110;
        rom_memory[6016] = 3'b110;
        rom_memory[6017] = 3'b110;
        rom_memory[6018] = 3'b110;
        rom_memory[6019] = 3'b110;
        rom_memory[6020] = 3'b110;
        rom_memory[6021] = 3'b110;
        rom_memory[6022] = 3'b110;
        rom_memory[6023] = 3'b110;
        rom_memory[6024] = 3'b110;
        rom_memory[6025] = 3'b110;
        rom_memory[6026] = 3'b110;
        rom_memory[6027] = 3'b110;
        rom_memory[6028] = 3'b110;
        rom_memory[6029] = 3'b110;
        rom_memory[6030] = 3'b110;
        rom_memory[6031] = 3'b110;
        rom_memory[6032] = 3'b000;
        rom_memory[6033] = 3'b000;
        rom_memory[6034] = 3'b000;
        rom_memory[6035] = 3'b000;
        rom_memory[6036] = 3'b000;
        rom_memory[6037] = 3'b000;
        rom_memory[6038] = 3'b000;
        rom_memory[6039] = 3'b000;
        rom_memory[6040] = 3'b111;
        rom_memory[6041] = 3'b111;
        rom_memory[6042] = 3'b111;
        rom_memory[6043] = 3'b111;
        rom_memory[6044] = 3'b111;
        rom_memory[6045] = 3'b111;
        rom_memory[6046] = 3'b111;
        rom_memory[6047] = 3'b111;
        rom_memory[6048] = 3'b110;
        rom_memory[6049] = 3'b110;
        rom_memory[6050] = 3'b111;
        rom_memory[6051] = 3'b111;
        rom_memory[6052] = 3'b111;
        rom_memory[6053] = 3'b111;
        rom_memory[6054] = 3'b111;
        rom_memory[6055] = 3'b000;
        rom_memory[6056] = 3'b000;
        rom_memory[6057] = 3'b000;
        rom_memory[6058] = 3'b000;
        rom_memory[6059] = 3'b000;
        rom_memory[6060] = 3'b000;
        rom_memory[6061] = 3'b000;
        rom_memory[6062] = 3'b000;
        rom_memory[6063] = 3'b000;
        rom_memory[6064] = 3'b000;
        rom_memory[6065] = 3'b000;
        rom_memory[6066] = 3'b000;
        rom_memory[6067] = 3'b000;
        rom_memory[6068] = 3'b000;
        rom_memory[6069] = 3'b000;
        rom_memory[6070] = 3'b000;
        rom_memory[6071] = 3'b000;
        rom_memory[6072] = 3'b000;
        rom_memory[6073] = 3'b011;
        rom_memory[6074] = 3'b000;
        rom_memory[6075] = 3'b001;
        rom_memory[6076] = 3'b011;
        rom_memory[6077] = 3'b011;
        rom_memory[6078] = 3'b011;
        rom_memory[6079] = 3'b011;
        rom_memory[6080] = 3'b011;
        rom_memory[6081] = 3'b011;
        rom_memory[6082] = 3'b111;
        rom_memory[6083] = 3'b111;
        rom_memory[6084] = 3'b111;
        rom_memory[6085] = 3'b110;
        rom_memory[6086] = 3'b110;
        rom_memory[6087] = 3'b110;
        rom_memory[6088] = 3'b110;
        rom_memory[6089] = 3'b110;
        rom_memory[6090] = 3'b110;
        rom_memory[6091] = 3'b110;
        rom_memory[6092] = 3'b110;
        rom_memory[6093] = 3'b110;
        rom_memory[6094] = 3'b110;
        rom_memory[6095] = 3'b110;
        rom_memory[6096] = 3'b110;
        rom_memory[6097] = 3'b110;
        rom_memory[6098] = 3'b110;
        rom_memory[6099] = 3'b110;
        rom_memory[6100] = 3'b110;
        rom_memory[6101] = 3'b110;
        rom_memory[6102] = 3'b110;
        rom_memory[6103] = 3'b110;
        rom_memory[6104] = 3'b110;
        rom_memory[6105] = 3'b110;
        rom_memory[6106] = 3'b110;
        rom_memory[6107] = 3'b110;
        rom_memory[6108] = 3'b110;
        rom_memory[6109] = 3'b110;
        rom_memory[6110] = 3'b110;
        rom_memory[6111] = 3'b110;
        rom_memory[6112] = 3'b110;
        rom_memory[6113] = 3'b110;
        rom_memory[6114] = 3'b110;
        rom_memory[6115] = 3'b110;
        rom_memory[6116] = 3'b110;
        rom_memory[6117] = 3'b110;
        rom_memory[6118] = 3'b110;
        rom_memory[6119] = 3'b110;
        rom_memory[6120] = 3'b110;
        rom_memory[6121] = 3'b110;
        rom_memory[6122] = 3'b110;
        rom_memory[6123] = 3'b110;
        rom_memory[6124] = 3'b110;
        rom_memory[6125] = 3'b110;
        rom_memory[6126] = 3'b110;
        rom_memory[6127] = 3'b110;
        rom_memory[6128] = 3'b110;
        rom_memory[6129] = 3'b110;
        rom_memory[6130] = 3'b110;
        rom_memory[6131] = 3'b110;
        rom_memory[6132] = 3'b110;
        rom_memory[6133] = 3'b110;
        rom_memory[6134] = 3'b110;
        rom_memory[6135] = 3'b110;
        rom_memory[6136] = 3'b110;
        rom_memory[6137] = 3'b110;
        rom_memory[6138] = 3'b110;
        rom_memory[6139] = 3'b110;
        rom_memory[6140] = 3'b110;
        rom_memory[6141] = 3'b110;
        rom_memory[6142] = 3'b110;
        rom_memory[6143] = 3'b110;
        rom_memory[6144] = 3'b110;
        rom_memory[6145] = 3'b110;
        rom_memory[6146] = 3'b110;
        rom_memory[6147] = 3'b110;
        rom_memory[6148] = 3'b110;
        rom_memory[6149] = 3'b110;
        rom_memory[6150] = 3'b110;
        rom_memory[6151] = 3'b110;
        rom_memory[6152] = 3'b110;
        rom_memory[6153] = 3'b110;
        rom_memory[6154] = 3'b110;
        rom_memory[6155] = 3'b110;
        rom_memory[6156] = 3'b110;
        rom_memory[6157] = 3'b110;
        rom_memory[6158] = 3'b110;
        rom_memory[6159] = 3'b110;
        rom_memory[6160] = 3'b110;
        rom_memory[6161] = 3'b110;
        rom_memory[6162] = 3'b110;
        rom_memory[6163] = 3'b110;
        rom_memory[6164] = 3'b110;
        rom_memory[6165] = 3'b110;
        rom_memory[6166] = 3'b110;
        rom_memory[6167] = 3'b110;
        rom_memory[6168] = 3'b110;
        rom_memory[6169] = 3'b110;
        rom_memory[6170] = 3'b110;
        rom_memory[6171] = 3'b110;
        rom_memory[6172] = 3'b110;
        rom_memory[6173] = 3'b110;
        rom_memory[6174] = 3'b110;
        rom_memory[6175] = 3'b110;
        rom_memory[6176] = 3'b110;
        rom_memory[6177] = 3'b110;
        rom_memory[6178] = 3'b110;
        rom_memory[6179] = 3'b110;
        rom_memory[6180] = 3'b110;
        rom_memory[6181] = 3'b110;
        rom_memory[6182] = 3'b110;
        rom_memory[6183] = 3'b110;
        rom_memory[6184] = 3'b110;
        rom_memory[6185] = 3'b110;
        rom_memory[6186] = 3'b110;
        rom_memory[6187] = 3'b110;
        rom_memory[6188] = 3'b110;
        rom_memory[6189] = 3'b110;
        rom_memory[6190] = 3'b110;
        rom_memory[6191] = 3'b110;
        rom_memory[6192] = 3'b110;
        rom_memory[6193] = 3'b110;
        rom_memory[6194] = 3'b110;
        rom_memory[6195] = 3'b110;
        rom_memory[6196] = 3'b110;
        rom_memory[6197] = 3'b110;
        rom_memory[6198] = 3'b110;
        rom_memory[6199] = 3'b110;
        rom_memory[6200] = 3'b110;
        rom_memory[6201] = 3'b110;
        rom_memory[6202] = 3'b110;
        rom_memory[6203] = 3'b110;
        rom_memory[6204] = 3'b110;
        rom_memory[6205] = 3'b110;
        rom_memory[6206] = 3'b110;
        rom_memory[6207] = 3'b110;
        rom_memory[6208] = 3'b110;
        rom_memory[6209] = 3'b110;
        rom_memory[6210] = 3'b110;
        rom_memory[6211] = 3'b110;
        rom_memory[6212] = 3'b110;
        rom_memory[6213] = 3'b110;
        rom_memory[6214] = 3'b110;
        rom_memory[6215] = 3'b110;
        rom_memory[6216] = 3'b110;
        rom_memory[6217] = 3'b110;
        rom_memory[6218] = 3'b110;
        rom_memory[6219] = 3'b110;
        rom_memory[6220] = 3'b110;
        rom_memory[6221] = 3'b110;
        rom_memory[6222] = 3'b110;
        rom_memory[6223] = 3'b110;
        rom_memory[6224] = 3'b110;
        rom_memory[6225] = 3'b110;
        rom_memory[6226] = 3'b110;
        rom_memory[6227] = 3'b110;
        rom_memory[6228] = 3'b110;
        rom_memory[6229] = 3'b110;
        rom_memory[6230] = 3'b110;
        rom_memory[6231] = 3'b110;
        rom_memory[6232] = 3'b110;
        rom_memory[6233] = 3'b110;
        rom_memory[6234] = 3'b110;
        rom_memory[6235] = 3'b110;
        rom_memory[6236] = 3'b110;
        rom_memory[6237] = 3'b110;
        rom_memory[6238] = 3'b110;
        rom_memory[6239] = 3'b110;
        rom_memory[6240] = 3'b110;
        rom_memory[6241] = 3'b110;
        rom_memory[6242] = 3'b110;
        rom_memory[6243] = 3'b110;
        rom_memory[6244] = 3'b110;
        rom_memory[6245] = 3'b110;
        rom_memory[6246] = 3'b110;
        rom_memory[6247] = 3'b110;
        rom_memory[6248] = 3'b110;
        rom_memory[6249] = 3'b110;
        rom_memory[6250] = 3'b110;
        rom_memory[6251] = 3'b110;
        rom_memory[6252] = 3'b110;
        rom_memory[6253] = 3'b110;
        rom_memory[6254] = 3'b110;
        rom_memory[6255] = 3'b110;
        rom_memory[6256] = 3'b110;
        rom_memory[6257] = 3'b110;
        rom_memory[6258] = 3'b110;
        rom_memory[6259] = 3'b110;
        rom_memory[6260] = 3'b110;
        rom_memory[6261] = 3'b110;
        rom_memory[6262] = 3'b110;
        rom_memory[6263] = 3'b110;
        rom_memory[6264] = 3'b110;
        rom_memory[6265] = 3'b110;
        rom_memory[6266] = 3'b110;
        rom_memory[6267] = 3'b110;
        rom_memory[6268] = 3'b110;
        rom_memory[6269] = 3'b110;
        rom_memory[6270] = 3'b110;
        rom_memory[6271] = 3'b110;
        rom_memory[6272] = 3'b110;
        rom_memory[6273] = 3'b110;
        rom_memory[6274] = 3'b100;
        rom_memory[6275] = 3'b000;
        rom_memory[6276] = 3'b000;
        rom_memory[6277] = 3'b000;
        rom_memory[6278] = 3'b000;
        rom_memory[6279] = 3'b000;
        rom_memory[6280] = 3'b000;
        rom_memory[6281] = 3'b111;
        rom_memory[6282] = 3'b111;
        rom_memory[6283] = 3'b111;
        rom_memory[6284] = 3'b111;
        rom_memory[6285] = 3'b111;
        rom_memory[6286] = 3'b111;
        rom_memory[6287] = 3'b111;
        rom_memory[6288] = 3'b111;
        rom_memory[6289] = 3'b111;
        rom_memory[6290] = 3'b111;
        rom_memory[6291] = 3'b111;
        rom_memory[6292] = 3'b111;
        rom_memory[6293] = 3'b111;
        rom_memory[6294] = 3'b111;
        rom_memory[6295] = 3'b000;
        rom_memory[6296] = 3'b000;
        rom_memory[6297] = 3'b000;
        rom_memory[6298] = 3'b000;
        rom_memory[6299] = 3'b000;
        rom_memory[6300] = 3'b000;
        rom_memory[6301] = 3'b000;
        rom_memory[6302] = 3'b000;
        rom_memory[6303] = 3'b000;
        rom_memory[6304] = 3'b000;
        rom_memory[6305] = 3'b000;
        rom_memory[6306] = 3'b000;
        rom_memory[6307] = 3'b000;
        rom_memory[6308] = 3'b000;
        rom_memory[6309] = 3'b000;
        rom_memory[6310] = 3'b000;
        rom_memory[6311] = 3'b000;
        rom_memory[6312] = 3'b000;
        rom_memory[6313] = 3'b000;
        rom_memory[6314] = 3'b000;
        rom_memory[6315] = 3'b011;
        rom_memory[6316] = 3'b000;
        rom_memory[6317] = 3'b011;
        rom_memory[6318] = 3'b011;
        rom_memory[6319] = 3'b011;
        rom_memory[6320] = 3'b011;
        rom_memory[6321] = 3'b011;
        rom_memory[6322] = 3'b011;
        rom_memory[6323] = 3'b111;
        rom_memory[6324] = 3'b111;
        rom_memory[6325] = 3'b111;
        rom_memory[6326] = 3'b110;
        rom_memory[6327] = 3'b110;
        rom_memory[6328] = 3'b110;
        rom_memory[6329] = 3'b110;
        rom_memory[6330] = 3'b110;
        rom_memory[6331] = 3'b110;
        rom_memory[6332] = 3'b110;
        rom_memory[6333] = 3'b110;
        rom_memory[6334] = 3'b110;
        rom_memory[6335] = 3'b110;
        rom_memory[6336] = 3'b110;
        rom_memory[6337] = 3'b110;
        rom_memory[6338] = 3'b110;
        rom_memory[6339] = 3'b110;
        rom_memory[6340] = 3'b110;
        rom_memory[6341] = 3'b110;
        rom_memory[6342] = 3'b110;
        rom_memory[6343] = 3'b110;
        rom_memory[6344] = 3'b110;
        rom_memory[6345] = 3'b110;
        rom_memory[6346] = 3'b110;
        rom_memory[6347] = 3'b110;
        rom_memory[6348] = 3'b110;
        rom_memory[6349] = 3'b110;
        rom_memory[6350] = 3'b110;
        rom_memory[6351] = 3'b110;
        rom_memory[6352] = 3'b110;
        rom_memory[6353] = 3'b110;
        rom_memory[6354] = 3'b110;
        rom_memory[6355] = 3'b110;
        rom_memory[6356] = 3'b110;
        rom_memory[6357] = 3'b110;
        rom_memory[6358] = 3'b110;
        rom_memory[6359] = 3'b110;
        rom_memory[6360] = 3'b110;
        rom_memory[6361] = 3'b110;
        rom_memory[6362] = 3'b110;
        rom_memory[6363] = 3'b110;
        rom_memory[6364] = 3'b110;
        rom_memory[6365] = 3'b110;
        rom_memory[6366] = 3'b110;
        rom_memory[6367] = 3'b110;
        rom_memory[6368] = 3'b110;
        rom_memory[6369] = 3'b110;
        rom_memory[6370] = 3'b110;
        rom_memory[6371] = 3'b110;
        rom_memory[6372] = 3'b110;
        rom_memory[6373] = 3'b110;
        rom_memory[6374] = 3'b110;
        rom_memory[6375] = 3'b110;
        rom_memory[6376] = 3'b110;
        rom_memory[6377] = 3'b110;
        rom_memory[6378] = 3'b110;
        rom_memory[6379] = 3'b110;
        rom_memory[6380] = 3'b110;
        rom_memory[6381] = 3'b110;
        rom_memory[6382] = 3'b110;
        rom_memory[6383] = 3'b110;
        rom_memory[6384] = 3'b110;
        rom_memory[6385] = 3'b110;
        rom_memory[6386] = 3'b110;
        rom_memory[6387] = 3'b110;
        rom_memory[6388] = 3'b110;
        rom_memory[6389] = 3'b110;
        rom_memory[6390] = 3'b110;
        rom_memory[6391] = 3'b110;
        rom_memory[6392] = 3'b110;
        rom_memory[6393] = 3'b110;
        rom_memory[6394] = 3'b110;
        rom_memory[6395] = 3'b110;
        rom_memory[6396] = 3'b110;
        rom_memory[6397] = 3'b110;
        rom_memory[6398] = 3'b110;
        rom_memory[6399] = 3'b110;
        rom_memory[6400] = 3'b110;
        rom_memory[6401] = 3'b110;
        rom_memory[6402] = 3'b110;
        rom_memory[6403] = 3'b110;
        rom_memory[6404] = 3'b110;
        rom_memory[6405] = 3'b110;
        rom_memory[6406] = 3'b110;
        rom_memory[6407] = 3'b110;
        rom_memory[6408] = 3'b110;
        rom_memory[6409] = 3'b110;
        rom_memory[6410] = 3'b110;
        rom_memory[6411] = 3'b110;
        rom_memory[6412] = 3'b110;
        rom_memory[6413] = 3'b110;
        rom_memory[6414] = 3'b110;
        rom_memory[6415] = 3'b110;
        rom_memory[6416] = 3'b110;
        rom_memory[6417] = 3'b110;
        rom_memory[6418] = 3'b110;
        rom_memory[6419] = 3'b110;
        rom_memory[6420] = 3'b110;
        rom_memory[6421] = 3'b110;
        rom_memory[6422] = 3'b110;
        rom_memory[6423] = 3'b110;
        rom_memory[6424] = 3'b110;
        rom_memory[6425] = 3'b110;
        rom_memory[6426] = 3'b110;
        rom_memory[6427] = 3'b110;
        rom_memory[6428] = 3'b110;
        rom_memory[6429] = 3'b110;
        rom_memory[6430] = 3'b110;
        rom_memory[6431] = 3'b110;
        rom_memory[6432] = 3'b110;
        rom_memory[6433] = 3'b110;
        rom_memory[6434] = 3'b110;
        rom_memory[6435] = 3'b110;
        rom_memory[6436] = 3'b110;
        rom_memory[6437] = 3'b110;
        rom_memory[6438] = 3'b110;
        rom_memory[6439] = 3'b110;
        rom_memory[6440] = 3'b110;
        rom_memory[6441] = 3'b110;
        rom_memory[6442] = 3'b110;
        rom_memory[6443] = 3'b110;
        rom_memory[6444] = 3'b110;
        rom_memory[6445] = 3'b110;
        rom_memory[6446] = 3'b110;
        rom_memory[6447] = 3'b110;
        rom_memory[6448] = 3'b110;
        rom_memory[6449] = 3'b110;
        rom_memory[6450] = 3'b110;
        rom_memory[6451] = 3'b110;
        rom_memory[6452] = 3'b110;
        rom_memory[6453] = 3'b110;
        rom_memory[6454] = 3'b110;
        rom_memory[6455] = 3'b110;
        rom_memory[6456] = 3'b110;
        rom_memory[6457] = 3'b110;
        rom_memory[6458] = 3'b110;
        rom_memory[6459] = 3'b110;
        rom_memory[6460] = 3'b110;
        rom_memory[6461] = 3'b110;
        rom_memory[6462] = 3'b110;
        rom_memory[6463] = 3'b110;
        rom_memory[6464] = 3'b110;
        rom_memory[6465] = 3'b110;
        rom_memory[6466] = 3'b110;
        rom_memory[6467] = 3'b110;
        rom_memory[6468] = 3'b110;
        rom_memory[6469] = 3'b110;
        rom_memory[6470] = 3'b110;
        rom_memory[6471] = 3'b110;
        rom_memory[6472] = 3'b110;
        rom_memory[6473] = 3'b110;
        rom_memory[6474] = 3'b110;
        rom_memory[6475] = 3'b110;
        rom_memory[6476] = 3'b110;
        rom_memory[6477] = 3'b110;
        rom_memory[6478] = 3'b110;
        rom_memory[6479] = 3'b110;
        rom_memory[6480] = 3'b110;
        rom_memory[6481] = 3'b110;
        rom_memory[6482] = 3'b110;
        rom_memory[6483] = 3'b110;
        rom_memory[6484] = 3'b110;
        rom_memory[6485] = 3'b110;
        rom_memory[6486] = 3'b110;
        rom_memory[6487] = 3'b110;
        rom_memory[6488] = 3'b110;
        rom_memory[6489] = 3'b110;
        rom_memory[6490] = 3'b110;
        rom_memory[6491] = 3'b110;
        rom_memory[6492] = 3'b110;
        rom_memory[6493] = 3'b110;
        rom_memory[6494] = 3'b110;
        rom_memory[6495] = 3'b110;
        rom_memory[6496] = 3'b110;
        rom_memory[6497] = 3'b110;
        rom_memory[6498] = 3'b110;
        rom_memory[6499] = 3'b110;
        rom_memory[6500] = 3'b110;
        rom_memory[6501] = 3'b110;
        rom_memory[6502] = 3'b110;
        rom_memory[6503] = 3'b110;
        rom_memory[6504] = 3'b110;
        rom_memory[6505] = 3'b110;
        rom_memory[6506] = 3'b110;
        rom_memory[6507] = 3'b110;
        rom_memory[6508] = 3'b110;
        rom_memory[6509] = 3'b110;
        rom_memory[6510] = 3'b110;
        rom_memory[6511] = 3'b110;
        rom_memory[6512] = 3'b110;
        rom_memory[6513] = 3'b110;
        rom_memory[6514] = 3'b110;
        rom_memory[6515] = 3'b110;
        rom_memory[6516] = 3'b110;
        rom_memory[6517] = 3'b000;
        rom_memory[6518] = 3'b000;
        rom_memory[6519] = 3'b000;
        rom_memory[6520] = 3'b000;
        rom_memory[6521] = 3'b000;
        rom_memory[6522] = 3'b000;
        rom_memory[6523] = 3'b111;
        rom_memory[6524] = 3'b111;
        rom_memory[6525] = 3'b111;
        rom_memory[6526] = 3'b111;
        rom_memory[6527] = 3'b111;
        rom_memory[6528] = 3'b111;
        rom_memory[6529] = 3'b111;
        rom_memory[6530] = 3'b111;
        rom_memory[6531] = 3'b111;
        rom_memory[6532] = 3'b111;
        rom_memory[6533] = 3'b111;
        rom_memory[6534] = 3'b111;
        rom_memory[6535] = 3'b000;
        rom_memory[6536] = 3'b000;
        rom_memory[6537] = 3'b000;
        rom_memory[6538] = 3'b000;
        rom_memory[6539] = 3'b000;
        rom_memory[6540] = 3'b000;
        rom_memory[6541] = 3'b000;
        rom_memory[6542] = 3'b000;
        rom_memory[6543] = 3'b000;
        rom_memory[6544] = 3'b000;
        rom_memory[6545] = 3'b000;
        rom_memory[6546] = 3'b000;
        rom_memory[6547] = 3'b000;
        rom_memory[6548] = 3'b000;
        rom_memory[6549] = 3'b000;
        rom_memory[6550] = 3'b000;
        rom_memory[6551] = 3'b000;
        rom_memory[6552] = 3'b000;
        rom_memory[6553] = 3'b000;
        rom_memory[6554] = 3'b010;
        rom_memory[6555] = 3'b000;
        rom_memory[6556] = 3'b000;
        rom_memory[6557] = 3'b011;
        rom_memory[6558] = 3'b011;
        rom_memory[6559] = 3'b011;
        rom_memory[6560] = 3'b011;
        rom_memory[6561] = 3'b011;
        rom_memory[6562] = 3'b011;
        rom_memory[6563] = 3'b111;
        rom_memory[6564] = 3'b111;
        rom_memory[6565] = 3'b111;
        rom_memory[6566] = 3'b111;
        rom_memory[6567] = 3'b110;
        rom_memory[6568] = 3'b110;
        rom_memory[6569] = 3'b110;
        rom_memory[6570] = 3'b110;
        rom_memory[6571] = 3'b110;
        rom_memory[6572] = 3'b110;
        rom_memory[6573] = 3'b110;
        rom_memory[6574] = 3'b110;
        rom_memory[6575] = 3'b110;
        rom_memory[6576] = 3'b110;
        rom_memory[6577] = 3'b110;
        rom_memory[6578] = 3'b110;
        rom_memory[6579] = 3'b110;
        rom_memory[6580] = 3'b110;
        rom_memory[6581] = 3'b110;
        rom_memory[6582] = 3'b110;
        rom_memory[6583] = 3'b110;
        rom_memory[6584] = 3'b110;
        rom_memory[6585] = 3'b110;
        rom_memory[6586] = 3'b110;
        rom_memory[6587] = 3'b110;
        rom_memory[6588] = 3'b110;
        rom_memory[6589] = 3'b110;
        rom_memory[6590] = 3'b110;
        rom_memory[6591] = 3'b110;
        rom_memory[6592] = 3'b110;
        rom_memory[6593] = 3'b110;
        rom_memory[6594] = 3'b110;
        rom_memory[6595] = 3'b110;
        rom_memory[6596] = 3'b110;
        rom_memory[6597] = 3'b110;
        rom_memory[6598] = 3'b110;
        rom_memory[6599] = 3'b110;
        rom_memory[6600] = 3'b110;
        rom_memory[6601] = 3'b110;
        rom_memory[6602] = 3'b110;
        rom_memory[6603] = 3'b110;
        rom_memory[6604] = 3'b110;
        rom_memory[6605] = 3'b110;
        rom_memory[6606] = 3'b110;
        rom_memory[6607] = 3'b110;
        rom_memory[6608] = 3'b110;
        rom_memory[6609] = 3'b110;
        rom_memory[6610] = 3'b110;
        rom_memory[6611] = 3'b110;
        rom_memory[6612] = 3'b110;
        rom_memory[6613] = 3'b110;
        rom_memory[6614] = 3'b110;
        rom_memory[6615] = 3'b110;
        rom_memory[6616] = 3'b110;
        rom_memory[6617] = 3'b110;
        rom_memory[6618] = 3'b110;
        rom_memory[6619] = 3'b110;
        rom_memory[6620] = 3'b110;
        rom_memory[6621] = 3'b110;
        rom_memory[6622] = 3'b110;
        rom_memory[6623] = 3'b110;
        rom_memory[6624] = 3'b110;
        rom_memory[6625] = 3'b110;
        rom_memory[6626] = 3'b110;
        rom_memory[6627] = 3'b110;
        rom_memory[6628] = 3'b110;
        rom_memory[6629] = 3'b110;
        rom_memory[6630] = 3'b110;
        rom_memory[6631] = 3'b110;
        rom_memory[6632] = 3'b110;
        rom_memory[6633] = 3'b110;
        rom_memory[6634] = 3'b110;
        rom_memory[6635] = 3'b110;
        rom_memory[6636] = 3'b110;
        rom_memory[6637] = 3'b110;
        rom_memory[6638] = 3'b110;
        rom_memory[6639] = 3'b110;
        rom_memory[6640] = 3'b110;
        rom_memory[6641] = 3'b110;
        rom_memory[6642] = 3'b110;
        rom_memory[6643] = 3'b110;
        rom_memory[6644] = 3'b110;
        rom_memory[6645] = 3'b110;
        rom_memory[6646] = 3'b110;
        rom_memory[6647] = 3'b110;
        rom_memory[6648] = 3'b110;
        rom_memory[6649] = 3'b110;
        rom_memory[6650] = 3'b110;
        rom_memory[6651] = 3'b110;
        rom_memory[6652] = 3'b110;
        rom_memory[6653] = 3'b110;
        rom_memory[6654] = 3'b110;
        rom_memory[6655] = 3'b110;
        rom_memory[6656] = 3'b110;
        rom_memory[6657] = 3'b110;
        rom_memory[6658] = 3'b110;
        rom_memory[6659] = 3'b110;
        rom_memory[6660] = 3'b110;
        rom_memory[6661] = 3'b110;
        rom_memory[6662] = 3'b110;
        rom_memory[6663] = 3'b110;
        rom_memory[6664] = 3'b110;
        rom_memory[6665] = 3'b110;
        rom_memory[6666] = 3'b110;
        rom_memory[6667] = 3'b110;
        rom_memory[6668] = 3'b110;
        rom_memory[6669] = 3'b110;
        rom_memory[6670] = 3'b110;
        rom_memory[6671] = 3'b110;
        rom_memory[6672] = 3'b110;
        rom_memory[6673] = 3'b110;
        rom_memory[6674] = 3'b110;
        rom_memory[6675] = 3'b110;
        rom_memory[6676] = 3'b110;
        rom_memory[6677] = 3'b110;
        rom_memory[6678] = 3'b110;
        rom_memory[6679] = 3'b110;
        rom_memory[6680] = 3'b110;
        rom_memory[6681] = 3'b110;
        rom_memory[6682] = 3'b110;
        rom_memory[6683] = 3'b110;
        rom_memory[6684] = 3'b110;
        rom_memory[6685] = 3'b110;
        rom_memory[6686] = 3'b110;
        rom_memory[6687] = 3'b110;
        rom_memory[6688] = 3'b110;
        rom_memory[6689] = 3'b110;
        rom_memory[6690] = 3'b110;
        rom_memory[6691] = 3'b110;
        rom_memory[6692] = 3'b110;
        rom_memory[6693] = 3'b110;
        rom_memory[6694] = 3'b110;
        rom_memory[6695] = 3'b110;
        rom_memory[6696] = 3'b110;
        rom_memory[6697] = 3'b110;
        rom_memory[6698] = 3'b110;
        rom_memory[6699] = 3'b110;
        rom_memory[6700] = 3'b110;
        rom_memory[6701] = 3'b110;
        rom_memory[6702] = 3'b110;
        rom_memory[6703] = 3'b110;
        rom_memory[6704] = 3'b110;
        rom_memory[6705] = 3'b110;
        rom_memory[6706] = 3'b110;
        rom_memory[6707] = 3'b110;
        rom_memory[6708] = 3'b110;
        rom_memory[6709] = 3'b110;
        rom_memory[6710] = 3'b110;
        rom_memory[6711] = 3'b110;
        rom_memory[6712] = 3'b110;
        rom_memory[6713] = 3'b110;
        rom_memory[6714] = 3'b110;
        rom_memory[6715] = 3'b110;
        rom_memory[6716] = 3'b110;
        rom_memory[6717] = 3'b110;
        rom_memory[6718] = 3'b110;
        rom_memory[6719] = 3'b110;
        rom_memory[6720] = 3'b110;
        rom_memory[6721] = 3'b110;
        rom_memory[6722] = 3'b110;
        rom_memory[6723] = 3'b110;
        rom_memory[6724] = 3'b110;
        rom_memory[6725] = 3'b110;
        rom_memory[6726] = 3'b110;
        rom_memory[6727] = 3'b110;
        rom_memory[6728] = 3'b110;
        rom_memory[6729] = 3'b110;
        rom_memory[6730] = 3'b110;
        rom_memory[6731] = 3'b110;
        rom_memory[6732] = 3'b110;
        rom_memory[6733] = 3'b110;
        rom_memory[6734] = 3'b110;
        rom_memory[6735] = 3'b110;
        rom_memory[6736] = 3'b110;
        rom_memory[6737] = 3'b110;
        rom_memory[6738] = 3'b110;
        rom_memory[6739] = 3'b110;
        rom_memory[6740] = 3'b110;
        rom_memory[6741] = 3'b110;
        rom_memory[6742] = 3'b110;
        rom_memory[6743] = 3'b110;
        rom_memory[6744] = 3'b110;
        rom_memory[6745] = 3'b110;
        rom_memory[6746] = 3'b110;
        rom_memory[6747] = 3'b110;
        rom_memory[6748] = 3'b110;
        rom_memory[6749] = 3'b110;
        rom_memory[6750] = 3'b110;
        rom_memory[6751] = 3'b110;
        rom_memory[6752] = 3'b110;
        rom_memory[6753] = 3'b110;
        rom_memory[6754] = 3'b110;
        rom_memory[6755] = 3'b110;
        rom_memory[6756] = 3'b110;
        rom_memory[6757] = 3'b110;
        rom_memory[6758] = 3'b110;
        rom_memory[6759] = 3'b000;
        rom_memory[6760] = 3'b000;
        rom_memory[6761] = 3'b000;
        rom_memory[6762] = 3'b000;
        rom_memory[6763] = 3'b000;
        rom_memory[6764] = 3'b101;
        rom_memory[6765] = 3'b111;
        rom_memory[6766] = 3'b000;
        rom_memory[6767] = 3'b000;
        rom_memory[6768] = 3'b111;
        rom_memory[6769] = 3'b111;
        rom_memory[6770] = 3'b111;
        rom_memory[6771] = 3'b111;
        rom_memory[6772] = 3'b111;
        rom_memory[6773] = 3'b111;
        rom_memory[6774] = 3'b000;
        rom_memory[6775] = 3'b000;
        rom_memory[6776] = 3'b000;
        rom_memory[6777] = 3'b000;
        rom_memory[6778] = 3'b000;
        rom_memory[6779] = 3'b000;
        rom_memory[6780] = 3'b000;
        rom_memory[6781] = 3'b000;
        rom_memory[6782] = 3'b000;
        rom_memory[6783] = 3'b000;
        rom_memory[6784] = 3'b000;
        rom_memory[6785] = 3'b000;
        rom_memory[6786] = 3'b000;
        rom_memory[6787] = 3'b000;
        rom_memory[6788] = 3'b000;
        rom_memory[6789] = 3'b000;
        rom_memory[6790] = 3'b000;
        rom_memory[6791] = 3'b000;
        rom_memory[6792] = 3'b000;
        rom_memory[6793] = 3'b000;
        rom_memory[6794] = 3'b010;
        rom_memory[6795] = 3'b000;
        rom_memory[6796] = 3'b011;
        rom_memory[6797] = 3'b011;
        rom_memory[6798] = 3'b011;
        rom_memory[6799] = 3'b011;
        rom_memory[6800] = 3'b010;
        rom_memory[6801] = 3'b000;
        rom_memory[6802] = 3'b011;
        rom_memory[6803] = 3'b011;
        rom_memory[6804] = 3'b111;
        rom_memory[6805] = 3'b111;
        rom_memory[6806] = 3'b111;
        rom_memory[6807] = 3'b111;
        rom_memory[6808] = 3'b111;
        rom_memory[6809] = 3'b110;
        rom_memory[6810] = 3'b110;
        rom_memory[6811] = 3'b110;
        rom_memory[6812] = 3'b110;
        rom_memory[6813] = 3'b110;
        rom_memory[6814] = 3'b110;
        rom_memory[6815] = 3'b110;
        rom_memory[6816] = 3'b110;
        rom_memory[6817] = 3'b110;
        rom_memory[6818] = 3'b110;
        rom_memory[6819] = 3'b110;
        rom_memory[6820] = 3'b110;
        rom_memory[6821] = 3'b110;
        rom_memory[6822] = 3'b110;
        rom_memory[6823] = 3'b110;
        rom_memory[6824] = 3'b110;
        rom_memory[6825] = 3'b110;
        rom_memory[6826] = 3'b110;
        rom_memory[6827] = 3'b110;
        rom_memory[6828] = 3'b110;
        rom_memory[6829] = 3'b110;
        rom_memory[6830] = 3'b110;
        rom_memory[6831] = 3'b110;
        rom_memory[6832] = 3'b110;
        rom_memory[6833] = 3'b110;
        rom_memory[6834] = 3'b110;
        rom_memory[6835] = 3'b110;
        rom_memory[6836] = 3'b110;
        rom_memory[6837] = 3'b110;
        rom_memory[6838] = 3'b110;
        rom_memory[6839] = 3'b110;
        rom_memory[6840] = 3'b110;
        rom_memory[6841] = 3'b110;
        rom_memory[6842] = 3'b110;
        rom_memory[6843] = 3'b110;
        rom_memory[6844] = 3'b110;
        rom_memory[6845] = 3'b110;
        rom_memory[6846] = 3'b110;
        rom_memory[6847] = 3'b110;
        rom_memory[6848] = 3'b110;
        rom_memory[6849] = 3'b110;
        rom_memory[6850] = 3'b110;
        rom_memory[6851] = 3'b110;
        rom_memory[6852] = 3'b110;
        rom_memory[6853] = 3'b110;
        rom_memory[6854] = 3'b110;
        rom_memory[6855] = 3'b110;
        rom_memory[6856] = 3'b110;
        rom_memory[6857] = 3'b110;
        rom_memory[6858] = 3'b110;
        rom_memory[6859] = 3'b110;
        rom_memory[6860] = 3'b110;
        rom_memory[6861] = 3'b110;
        rom_memory[6862] = 3'b110;
        rom_memory[6863] = 3'b110;
        rom_memory[6864] = 3'b110;
        rom_memory[6865] = 3'b110;
        rom_memory[6866] = 3'b110;
        rom_memory[6867] = 3'b110;
        rom_memory[6868] = 3'b110;
        rom_memory[6869] = 3'b110;
        rom_memory[6870] = 3'b110;
        rom_memory[6871] = 3'b110;
        rom_memory[6872] = 3'b110;
        rom_memory[6873] = 3'b110;
        rom_memory[6874] = 3'b110;
        rom_memory[6875] = 3'b110;
        rom_memory[6876] = 3'b110;
        rom_memory[6877] = 3'b110;
        rom_memory[6878] = 3'b110;
        rom_memory[6879] = 3'b110;
        rom_memory[6880] = 3'b110;
        rom_memory[6881] = 3'b110;
        rom_memory[6882] = 3'b110;
        rom_memory[6883] = 3'b110;
        rom_memory[6884] = 3'b110;
        rom_memory[6885] = 3'b110;
        rom_memory[6886] = 3'b110;
        rom_memory[6887] = 3'b110;
        rom_memory[6888] = 3'b110;
        rom_memory[6889] = 3'b110;
        rom_memory[6890] = 3'b110;
        rom_memory[6891] = 3'b110;
        rom_memory[6892] = 3'b110;
        rom_memory[6893] = 3'b110;
        rom_memory[6894] = 3'b110;
        rom_memory[6895] = 3'b110;
        rom_memory[6896] = 3'b110;
        rom_memory[6897] = 3'b110;
        rom_memory[6898] = 3'b110;
        rom_memory[6899] = 3'b110;
        rom_memory[6900] = 3'b110;
        rom_memory[6901] = 3'b110;
        rom_memory[6902] = 3'b110;
        rom_memory[6903] = 3'b110;
        rom_memory[6904] = 3'b110;
        rom_memory[6905] = 3'b110;
        rom_memory[6906] = 3'b110;
        rom_memory[6907] = 3'b110;
        rom_memory[6908] = 3'b110;
        rom_memory[6909] = 3'b110;
        rom_memory[6910] = 3'b110;
        rom_memory[6911] = 3'b110;
        rom_memory[6912] = 3'b110;
        rom_memory[6913] = 3'b110;
        rom_memory[6914] = 3'b110;
        rom_memory[6915] = 3'b110;
        rom_memory[6916] = 3'b110;
        rom_memory[6917] = 3'b110;
        rom_memory[6918] = 3'b110;
        rom_memory[6919] = 3'b110;
        rom_memory[6920] = 3'b110;
        rom_memory[6921] = 3'b110;
        rom_memory[6922] = 3'b110;
        rom_memory[6923] = 3'b110;
        rom_memory[6924] = 3'b110;
        rom_memory[6925] = 3'b110;
        rom_memory[6926] = 3'b110;
        rom_memory[6927] = 3'b110;
        rom_memory[6928] = 3'b110;
        rom_memory[6929] = 3'b110;
        rom_memory[6930] = 3'b110;
        rom_memory[6931] = 3'b110;
        rom_memory[6932] = 3'b110;
        rom_memory[6933] = 3'b110;
        rom_memory[6934] = 3'b110;
        rom_memory[6935] = 3'b110;
        rom_memory[6936] = 3'b110;
        rom_memory[6937] = 3'b110;
        rom_memory[6938] = 3'b110;
        rom_memory[6939] = 3'b110;
        rom_memory[6940] = 3'b110;
        rom_memory[6941] = 3'b110;
        rom_memory[6942] = 3'b110;
        rom_memory[6943] = 3'b110;
        rom_memory[6944] = 3'b110;
        rom_memory[6945] = 3'b110;
        rom_memory[6946] = 3'b110;
        rom_memory[6947] = 3'b110;
        rom_memory[6948] = 3'b110;
        rom_memory[6949] = 3'b110;
        rom_memory[6950] = 3'b110;
        rom_memory[6951] = 3'b110;
        rom_memory[6952] = 3'b110;
        rom_memory[6953] = 3'b110;
        rom_memory[6954] = 3'b110;
        rom_memory[6955] = 3'b110;
        rom_memory[6956] = 3'b110;
        rom_memory[6957] = 3'b110;
        rom_memory[6958] = 3'b110;
        rom_memory[6959] = 3'b110;
        rom_memory[6960] = 3'b110;
        rom_memory[6961] = 3'b110;
        rom_memory[6962] = 3'b110;
        rom_memory[6963] = 3'b110;
        rom_memory[6964] = 3'b110;
        rom_memory[6965] = 3'b110;
        rom_memory[6966] = 3'b110;
        rom_memory[6967] = 3'b110;
        rom_memory[6968] = 3'b110;
        rom_memory[6969] = 3'b110;
        rom_memory[6970] = 3'b110;
        rom_memory[6971] = 3'b110;
        rom_memory[6972] = 3'b110;
        rom_memory[6973] = 3'b110;
        rom_memory[6974] = 3'b110;
        rom_memory[6975] = 3'b110;
        rom_memory[6976] = 3'b110;
        rom_memory[6977] = 3'b110;
        rom_memory[6978] = 3'b110;
        rom_memory[6979] = 3'b110;
        rom_memory[6980] = 3'b110;
        rom_memory[6981] = 3'b110;
        rom_memory[6982] = 3'b110;
        rom_memory[6983] = 3'b110;
        rom_memory[6984] = 3'b110;
        rom_memory[6985] = 3'b110;
        rom_memory[6986] = 3'b110;
        rom_memory[6987] = 3'b110;
        rom_memory[6988] = 3'b110;
        rom_memory[6989] = 3'b110;
        rom_memory[6990] = 3'b110;
        rom_memory[6991] = 3'b110;
        rom_memory[6992] = 3'b110;
        rom_memory[6993] = 3'b110;
        rom_memory[6994] = 3'b110;
        rom_memory[6995] = 3'b110;
        rom_memory[6996] = 3'b110;
        rom_memory[6997] = 3'b110;
        rom_memory[6998] = 3'b110;
        rom_memory[6999] = 3'b110;
        rom_memory[7000] = 3'b110;
        rom_memory[7001] = 3'b000;
        rom_memory[7002] = 3'b000;
        rom_memory[7003] = 3'b000;
        rom_memory[7004] = 3'b000;
        rom_memory[7005] = 3'b000;
        rom_memory[7006] = 3'b111;
        rom_memory[7007] = 3'b111;
        rom_memory[7008] = 3'b000;
        rom_memory[7009] = 3'b000;
        rom_memory[7010] = 3'b000;
        rom_memory[7011] = 3'b111;
        rom_memory[7012] = 3'b111;
        rom_memory[7013] = 3'b111;
        rom_memory[7014] = 3'b000;
        rom_memory[7015] = 3'b000;
        rom_memory[7016] = 3'b000;
        rom_memory[7017] = 3'b000;
        rom_memory[7018] = 3'b000;
        rom_memory[7019] = 3'b000;
        rom_memory[7020] = 3'b000;
        rom_memory[7021] = 3'b000;
        rom_memory[7022] = 3'b000;
        rom_memory[7023] = 3'b000;
        rom_memory[7024] = 3'b000;
        rom_memory[7025] = 3'b000;
        rom_memory[7026] = 3'b000;
        rom_memory[7027] = 3'b000;
        rom_memory[7028] = 3'b000;
        rom_memory[7029] = 3'b000;
        rom_memory[7030] = 3'b000;
        rom_memory[7031] = 3'b000;
        rom_memory[7032] = 3'b000;
        rom_memory[7033] = 3'b000;
        rom_memory[7034] = 3'b010;
        rom_memory[7035] = 3'b000;
        rom_memory[7036] = 3'b011;
        rom_memory[7037] = 3'b011;
        rom_memory[7038] = 3'b011;
        rom_memory[7039] = 3'b011;
        rom_memory[7040] = 3'b011;
        rom_memory[7041] = 3'b011;
        rom_memory[7042] = 3'b011;
        rom_memory[7043] = 3'b011;
        rom_memory[7044] = 3'b011;
        rom_memory[7045] = 3'b011;
        rom_memory[7046] = 3'b111;
        rom_memory[7047] = 3'b111;
        rom_memory[7048] = 3'b111;
        rom_memory[7049] = 3'b111;
        rom_memory[7050] = 3'b110;
        rom_memory[7051] = 3'b111;
        rom_memory[7052] = 3'b110;
        rom_memory[7053] = 3'b110;
        rom_memory[7054] = 3'b110;
        rom_memory[7055] = 3'b110;
        rom_memory[7056] = 3'b110;
        rom_memory[7057] = 3'b110;
        rom_memory[7058] = 3'b110;
        rom_memory[7059] = 3'b110;
        rom_memory[7060] = 3'b110;
        rom_memory[7061] = 3'b110;
        rom_memory[7062] = 3'b110;
        rom_memory[7063] = 3'b110;
        rom_memory[7064] = 3'b110;
        rom_memory[7065] = 3'b110;
        rom_memory[7066] = 3'b110;
        rom_memory[7067] = 3'b110;
        rom_memory[7068] = 3'b110;
        rom_memory[7069] = 3'b110;
        rom_memory[7070] = 3'b110;
        rom_memory[7071] = 3'b110;
        rom_memory[7072] = 3'b110;
        rom_memory[7073] = 3'b110;
        rom_memory[7074] = 3'b110;
        rom_memory[7075] = 3'b110;
        rom_memory[7076] = 3'b110;
        rom_memory[7077] = 3'b110;
        rom_memory[7078] = 3'b110;
        rom_memory[7079] = 3'b110;
        rom_memory[7080] = 3'b110;
        rom_memory[7081] = 3'b110;
        rom_memory[7082] = 3'b110;
        rom_memory[7083] = 3'b110;
        rom_memory[7084] = 3'b110;
        rom_memory[7085] = 3'b110;
        rom_memory[7086] = 3'b110;
        rom_memory[7087] = 3'b110;
        rom_memory[7088] = 3'b110;
        rom_memory[7089] = 3'b110;
        rom_memory[7090] = 3'b110;
        rom_memory[7091] = 3'b110;
        rom_memory[7092] = 3'b110;
        rom_memory[7093] = 3'b110;
        rom_memory[7094] = 3'b110;
        rom_memory[7095] = 3'b110;
        rom_memory[7096] = 3'b110;
        rom_memory[7097] = 3'b110;
        rom_memory[7098] = 3'b110;
        rom_memory[7099] = 3'b110;
        rom_memory[7100] = 3'b110;
        rom_memory[7101] = 3'b110;
        rom_memory[7102] = 3'b110;
        rom_memory[7103] = 3'b110;
        rom_memory[7104] = 3'b110;
        rom_memory[7105] = 3'b110;
        rom_memory[7106] = 3'b110;
        rom_memory[7107] = 3'b110;
        rom_memory[7108] = 3'b110;
        rom_memory[7109] = 3'b110;
        rom_memory[7110] = 3'b110;
        rom_memory[7111] = 3'b110;
        rom_memory[7112] = 3'b110;
        rom_memory[7113] = 3'b110;
        rom_memory[7114] = 3'b110;
        rom_memory[7115] = 3'b110;
        rom_memory[7116] = 3'b110;
        rom_memory[7117] = 3'b110;
        rom_memory[7118] = 3'b110;
        rom_memory[7119] = 3'b110;
        rom_memory[7120] = 3'b110;
        rom_memory[7121] = 3'b110;
        rom_memory[7122] = 3'b110;
        rom_memory[7123] = 3'b110;
        rom_memory[7124] = 3'b110;
        rom_memory[7125] = 3'b110;
        rom_memory[7126] = 3'b110;
        rom_memory[7127] = 3'b110;
        rom_memory[7128] = 3'b110;
        rom_memory[7129] = 3'b110;
        rom_memory[7130] = 3'b110;
        rom_memory[7131] = 3'b110;
        rom_memory[7132] = 3'b110;
        rom_memory[7133] = 3'b110;
        rom_memory[7134] = 3'b110;
        rom_memory[7135] = 3'b110;
        rom_memory[7136] = 3'b110;
        rom_memory[7137] = 3'b110;
        rom_memory[7138] = 3'b110;
        rom_memory[7139] = 3'b110;
        rom_memory[7140] = 3'b110;
        rom_memory[7141] = 3'b110;
        rom_memory[7142] = 3'b110;
        rom_memory[7143] = 3'b110;
        rom_memory[7144] = 3'b110;
        rom_memory[7145] = 3'b110;
        rom_memory[7146] = 3'b110;
        rom_memory[7147] = 3'b110;
        rom_memory[7148] = 3'b110;
        rom_memory[7149] = 3'b110;
        rom_memory[7150] = 3'b110;
        rom_memory[7151] = 3'b110;
        rom_memory[7152] = 3'b110;
        rom_memory[7153] = 3'b110;
        rom_memory[7154] = 3'b110;
        rom_memory[7155] = 3'b110;
        rom_memory[7156] = 3'b110;
        rom_memory[7157] = 3'b110;
        rom_memory[7158] = 3'b110;
        rom_memory[7159] = 3'b110;
        rom_memory[7160] = 3'b110;
        rom_memory[7161] = 3'b110;
        rom_memory[7162] = 3'b110;
        rom_memory[7163] = 3'b110;
        rom_memory[7164] = 3'b110;
        rom_memory[7165] = 3'b110;
        rom_memory[7166] = 3'b110;
        rom_memory[7167] = 3'b110;
        rom_memory[7168] = 3'b110;
        rom_memory[7169] = 3'b110;
        rom_memory[7170] = 3'b110;
        rom_memory[7171] = 3'b110;
        rom_memory[7172] = 3'b110;
        rom_memory[7173] = 3'b110;
        rom_memory[7174] = 3'b110;
        rom_memory[7175] = 3'b110;
        rom_memory[7176] = 3'b110;
        rom_memory[7177] = 3'b110;
        rom_memory[7178] = 3'b110;
        rom_memory[7179] = 3'b110;
        rom_memory[7180] = 3'b110;
        rom_memory[7181] = 3'b110;
        rom_memory[7182] = 3'b110;
        rom_memory[7183] = 3'b110;
        rom_memory[7184] = 3'b110;
        rom_memory[7185] = 3'b110;
        rom_memory[7186] = 3'b110;
        rom_memory[7187] = 3'b110;
        rom_memory[7188] = 3'b110;
        rom_memory[7189] = 3'b110;
        rom_memory[7190] = 3'b110;
        rom_memory[7191] = 3'b110;
        rom_memory[7192] = 3'b110;
        rom_memory[7193] = 3'b110;
        rom_memory[7194] = 3'b110;
        rom_memory[7195] = 3'b110;
        rom_memory[7196] = 3'b110;
        rom_memory[7197] = 3'b110;
        rom_memory[7198] = 3'b110;
        rom_memory[7199] = 3'b110;
        rom_memory[7200] = 3'b110;
        rom_memory[7201] = 3'b110;
        rom_memory[7202] = 3'b110;
        rom_memory[7203] = 3'b110;
        rom_memory[7204] = 3'b110;
        rom_memory[7205] = 3'b110;
        rom_memory[7206] = 3'b110;
        rom_memory[7207] = 3'b110;
        rom_memory[7208] = 3'b110;
        rom_memory[7209] = 3'b110;
        rom_memory[7210] = 3'b110;
        rom_memory[7211] = 3'b110;
        rom_memory[7212] = 3'b110;
        rom_memory[7213] = 3'b110;
        rom_memory[7214] = 3'b110;
        rom_memory[7215] = 3'b110;
        rom_memory[7216] = 3'b110;
        rom_memory[7217] = 3'b110;
        rom_memory[7218] = 3'b110;
        rom_memory[7219] = 3'b110;
        rom_memory[7220] = 3'b110;
        rom_memory[7221] = 3'b110;
        rom_memory[7222] = 3'b110;
        rom_memory[7223] = 3'b110;
        rom_memory[7224] = 3'b110;
        rom_memory[7225] = 3'b110;
        rom_memory[7226] = 3'b110;
        rom_memory[7227] = 3'b110;
        rom_memory[7228] = 3'b110;
        rom_memory[7229] = 3'b110;
        rom_memory[7230] = 3'b110;
        rom_memory[7231] = 3'b110;
        rom_memory[7232] = 3'b110;
        rom_memory[7233] = 3'b110;
        rom_memory[7234] = 3'b110;
        rom_memory[7235] = 3'b110;
        rom_memory[7236] = 3'b110;
        rom_memory[7237] = 3'b110;
        rom_memory[7238] = 3'b110;
        rom_memory[7239] = 3'b110;
        rom_memory[7240] = 3'b110;
        rom_memory[7241] = 3'b110;
        rom_memory[7242] = 3'b100;
        rom_memory[7243] = 3'b000;
        rom_memory[7244] = 3'b000;
        rom_memory[7245] = 3'b000;
        rom_memory[7246] = 3'b000;
        rom_memory[7247] = 3'b111;
        rom_memory[7248] = 3'b111;
        rom_memory[7249] = 3'b111;
        rom_memory[7250] = 3'b111;
        rom_memory[7251] = 3'b000;
        rom_memory[7252] = 3'b000;
        rom_memory[7253] = 3'b000;
        rom_memory[7254] = 3'b000;
        rom_memory[7255] = 3'b000;
        rom_memory[7256] = 3'b000;
        rom_memory[7257] = 3'b000;
        rom_memory[7258] = 3'b000;
        rom_memory[7259] = 3'b000;
        rom_memory[7260] = 3'b000;
        rom_memory[7261] = 3'b000;
        rom_memory[7262] = 3'b000;
        rom_memory[7263] = 3'b000;
        rom_memory[7264] = 3'b000;
        rom_memory[7265] = 3'b000;
        rom_memory[7266] = 3'b000;
        rom_memory[7267] = 3'b000;
        rom_memory[7268] = 3'b000;
        rom_memory[7269] = 3'b000;
        rom_memory[7270] = 3'b000;
        rom_memory[7271] = 3'b000;
        rom_memory[7272] = 3'b000;
        rom_memory[7273] = 3'b000;
        rom_memory[7274] = 3'b000;
        rom_memory[7275] = 3'b000;
        rom_memory[7276] = 3'b011;
        rom_memory[7277] = 3'b000;
        rom_memory[7278] = 3'b011;
        rom_memory[7279] = 3'b010;
        rom_memory[7280] = 3'b010;
        rom_memory[7281] = 3'b011;
        rom_memory[7282] = 3'b011;
        rom_memory[7283] = 3'b011;
        rom_memory[7284] = 3'b011;
        rom_memory[7285] = 3'b011;
        rom_memory[7286] = 3'b011;
        rom_memory[7287] = 3'b111;
        rom_memory[7288] = 3'b111;
        rom_memory[7289] = 3'b111;
        rom_memory[7290] = 3'b111;
        rom_memory[7291] = 3'b110;
        rom_memory[7292] = 3'b110;
        rom_memory[7293] = 3'b110;
        rom_memory[7294] = 3'b110;
        rom_memory[7295] = 3'b110;
        rom_memory[7296] = 3'b110;
        rom_memory[7297] = 3'b110;
        rom_memory[7298] = 3'b110;
        rom_memory[7299] = 3'b110;
        rom_memory[7300] = 3'b110;
        rom_memory[7301] = 3'b110;
        rom_memory[7302] = 3'b110;
        rom_memory[7303] = 3'b110;
        rom_memory[7304] = 3'b110;
        rom_memory[7305] = 3'b110;
        rom_memory[7306] = 3'b110;
        rom_memory[7307] = 3'b110;
        rom_memory[7308] = 3'b110;
        rom_memory[7309] = 3'b110;
        rom_memory[7310] = 3'b110;
        rom_memory[7311] = 3'b110;
        rom_memory[7312] = 3'b110;
        rom_memory[7313] = 3'b110;
        rom_memory[7314] = 3'b110;
        rom_memory[7315] = 3'b110;
        rom_memory[7316] = 3'b110;
        rom_memory[7317] = 3'b110;
        rom_memory[7318] = 3'b110;
        rom_memory[7319] = 3'b110;
        rom_memory[7320] = 3'b110;
        rom_memory[7321] = 3'b110;
        rom_memory[7322] = 3'b110;
        rom_memory[7323] = 3'b110;
        rom_memory[7324] = 3'b110;
        rom_memory[7325] = 3'b110;
        rom_memory[7326] = 3'b110;
        rom_memory[7327] = 3'b110;
        rom_memory[7328] = 3'b110;
        rom_memory[7329] = 3'b110;
        rom_memory[7330] = 3'b110;
        rom_memory[7331] = 3'b110;
        rom_memory[7332] = 3'b110;
        rom_memory[7333] = 3'b110;
        rom_memory[7334] = 3'b110;
        rom_memory[7335] = 3'b110;
        rom_memory[7336] = 3'b110;
        rom_memory[7337] = 3'b110;
        rom_memory[7338] = 3'b110;
        rom_memory[7339] = 3'b110;
        rom_memory[7340] = 3'b110;
        rom_memory[7341] = 3'b110;
        rom_memory[7342] = 3'b110;
        rom_memory[7343] = 3'b110;
        rom_memory[7344] = 3'b110;
        rom_memory[7345] = 3'b110;
        rom_memory[7346] = 3'b110;
        rom_memory[7347] = 3'b110;
        rom_memory[7348] = 3'b110;
        rom_memory[7349] = 3'b110;
        rom_memory[7350] = 3'b110;
        rom_memory[7351] = 3'b110;
        rom_memory[7352] = 3'b110;
        rom_memory[7353] = 3'b110;
        rom_memory[7354] = 3'b110;
        rom_memory[7355] = 3'b110;
        rom_memory[7356] = 3'b110;
        rom_memory[7357] = 3'b110;
        rom_memory[7358] = 3'b110;
        rom_memory[7359] = 3'b110;
        rom_memory[7360] = 3'b110;
        rom_memory[7361] = 3'b110;
        rom_memory[7362] = 3'b110;
        rom_memory[7363] = 3'b110;
        rom_memory[7364] = 3'b110;
        rom_memory[7365] = 3'b110;
        rom_memory[7366] = 3'b110;
        rom_memory[7367] = 3'b110;
        rom_memory[7368] = 3'b110;
        rom_memory[7369] = 3'b110;
        rom_memory[7370] = 3'b110;
        rom_memory[7371] = 3'b110;
        rom_memory[7372] = 3'b110;
        rom_memory[7373] = 3'b110;
        rom_memory[7374] = 3'b110;
        rom_memory[7375] = 3'b110;
        rom_memory[7376] = 3'b110;
        rom_memory[7377] = 3'b110;
        rom_memory[7378] = 3'b110;
        rom_memory[7379] = 3'b110;
        rom_memory[7380] = 3'b110;
        rom_memory[7381] = 3'b110;
        rom_memory[7382] = 3'b110;
        rom_memory[7383] = 3'b110;
        rom_memory[7384] = 3'b110;
        rom_memory[7385] = 3'b110;
        rom_memory[7386] = 3'b110;
        rom_memory[7387] = 3'b110;
        rom_memory[7388] = 3'b110;
        rom_memory[7389] = 3'b110;
        rom_memory[7390] = 3'b110;
        rom_memory[7391] = 3'b110;
        rom_memory[7392] = 3'b110;
        rom_memory[7393] = 3'b110;
        rom_memory[7394] = 3'b110;
        rom_memory[7395] = 3'b110;
        rom_memory[7396] = 3'b110;
        rom_memory[7397] = 3'b110;
        rom_memory[7398] = 3'b110;
        rom_memory[7399] = 3'b110;
        rom_memory[7400] = 3'b110;
        rom_memory[7401] = 3'b110;
        rom_memory[7402] = 3'b110;
        rom_memory[7403] = 3'b110;
        rom_memory[7404] = 3'b110;
        rom_memory[7405] = 3'b110;
        rom_memory[7406] = 3'b110;
        rom_memory[7407] = 3'b110;
        rom_memory[7408] = 3'b110;
        rom_memory[7409] = 3'b110;
        rom_memory[7410] = 3'b110;
        rom_memory[7411] = 3'b110;
        rom_memory[7412] = 3'b110;
        rom_memory[7413] = 3'b110;
        rom_memory[7414] = 3'b110;
        rom_memory[7415] = 3'b110;
        rom_memory[7416] = 3'b110;
        rom_memory[7417] = 3'b110;
        rom_memory[7418] = 3'b110;
        rom_memory[7419] = 3'b110;
        rom_memory[7420] = 3'b110;
        rom_memory[7421] = 3'b110;
        rom_memory[7422] = 3'b110;
        rom_memory[7423] = 3'b110;
        rom_memory[7424] = 3'b110;
        rom_memory[7425] = 3'b110;
        rom_memory[7426] = 3'b110;
        rom_memory[7427] = 3'b110;
        rom_memory[7428] = 3'b110;
        rom_memory[7429] = 3'b110;
        rom_memory[7430] = 3'b110;
        rom_memory[7431] = 3'b110;
        rom_memory[7432] = 3'b110;
        rom_memory[7433] = 3'b110;
        rom_memory[7434] = 3'b110;
        rom_memory[7435] = 3'b110;
        rom_memory[7436] = 3'b110;
        rom_memory[7437] = 3'b110;
        rom_memory[7438] = 3'b110;
        rom_memory[7439] = 3'b110;
        rom_memory[7440] = 3'b110;
        rom_memory[7441] = 3'b110;
        rom_memory[7442] = 3'b110;
        rom_memory[7443] = 3'b110;
        rom_memory[7444] = 3'b110;
        rom_memory[7445] = 3'b110;
        rom_memory[7446] = 3'b110;
        rom_memory[7447] = 3'b110;
        rom_memory[7448] = 3'b110;
        rom_memory[7449] = 3'b110;
        rom_memory[7450] = 3'b110;
        rom_memory[7451] = 3'b110;
        rom_memory[7452] = 3'b110;
        rom_memory[7453] = 3'b110;
        rom_memory[7454] = 3'b110;
        rom_memory[7455] = 3'b110;
        rom_memory[7456] = 3'b110;
        rom_memory[7457] = 3'b110;
        rom_memory[7458] = 3'b110;
        rom_memory[7459] = 3'b110;
        rom_memory[7460] = 3'b110;
        rom_memory[7461] = 3'b110;
        rom_memory[7462] = 3'b110;
        rom_memory[7463] = 3'b110;
        rom_memory[7464] = 3'b110;
        rom_memory[7465] = 3'b110;
        rom_memory[7466] = 3'b110;
        rom_memory[7467] = 3'b110;
        rom_memory[7468] = 3'b110;
        rom_memory[7469] = 3'b110;
        rom_memory[7470] = 3'b110;
        rom_memory[7471] = 3'b110;
        rom_memory[7472] = 3'b110;
        rom_memory[7473] = 3'b110;
        rom_memory[7474] = 3'b110;
        rom_memory[7475] = 3'b110;
        rom_memory[7476] = 3'b110;
        rom_memory[7477] = 3'b110;
        rom_memory[7478] = 3'b110;
        rom_memory[7479] = 3'b110;
        rom_memory[7480] = 3'b110;
        rom_memory[7481] = 3'b110;
        rom_memory[7482] = 3'b110;
        rom_memory[7483] = 3'b110;
        rom_memory[7484] = 3'b000;
        rom_memory[7485] = 3'b000;
        rom_memory[7486] = 3'b000;
        rom_memory[7487] = 3'b000;
        rom_memory[7488] = 3'b111;
        rom_memory[7489] = 3'b111;
        rom_memory[7490] = 3'b111;
        rom_memory[7491] = 3'b000;
        rom_memory[7492] = 3'b000;
        rom_memory[7493] = 3'b000;
        rom_memory[7494] = 3'b000;
        rom_memory[7495] = 3'b000;
        rom_memory[7496] = 3'b000;
        rom_memory[7497] = 3'b000;
        rom_memory[7498] = 3'b000;
        rom_memory[7499] = 3'b000;
        rom_memory[7500] = 3'b000;
        rom_memory[7501] = 3'b000;
        rom_memory[7502] = 3'b000;
        rom_memory[7503] = 3'b000;
        rom_memory[7504] = 3'b000;
        rom_memory[7505] = 3'b000;
        rom_memory[7506] = 3'b000;
        rom_memory[7507] = 3'b000;
        rom_memory[7508] = 3'b000;
        rom_memory[7509] = 3'b000;
        rom_memory[7510] = 3'b000;
        rom_memory[7511] = 3'b000;
        rom_memory[7512] = 3'b000;
        rom_memory[7513] = 3'b000;
        rom_memory[7514] = 3'b000;
        rom_memory[7515] = 3'b000;
        rom_memory[7516] = 3'b000;
        rom_memory[7517] = 3'b000;
        rom_memory[7518] = 3'b010;
        rom_memory[7519] = 3'b000;
        rom_memory[7520] = 3'b010;
        rom_memory[7521] = 3'b010;
        rom_memory[7522] = 3'b011;
        rom_memory[7523] = 3'b011;
        rom_memory[7524] = 3'b011;
        rom_memory[7525] = 3'b011;
        rom_memory[7526] = 3'b001;
        rom_memory[7527] = 3'b011;
        rom_memory[7528] = 3'b011;
        rom_memory[7529] = 3'b111;
        rom_memory[7530] = 3'b111;
        rom_memory[7531] = 3'b111;
        rom_memory[7532] = 3'b110;
        rom_memory[7533] = 3'b110;
        rom_memory[7534] = 3'b110;
        rom_memory[7535] = 3'b110;
        rom_memory[7536] = 3'b110;
        rom_memory[7537] = 3'b110;
        rom_memory[7538] = 3'b110;
        rom_memory[7539] = 3'b110;
        rom_memory[7540] = 3'b110;
        rom_memory[7541] = 3'b110;
        rom_memory[7542] = 3'b110;
        rom_memory[7543] = 3'b110;
        rom_memory[7544] = 3'b110;
        rom_memory[7545] = 3'b110;
        rom_memory[7546] = 3'b110;
        rom_memory[7547] = 3'b110;
        rom_memory[7548] = 3'b110;
        rom_memory[7549] = 3'b110;
        rom_memory[7550] = 3'b110;
        rom_memory[7551] = 3'b110;
        rom_memory[7552] = 3'b110;
        rom_memory[7553] = 3'b110;
        rom_memory[7554] = 3'b110;
        rom_memory[7555] = 3'b110;
        rom_memory[7556] = 3'b110;
        rom_memory[7557] = 3'b110;
        rom_memory[7558] = 3'b110;
        rom_memory[7559] = 3'b110;
        rom_memory[7560] = 3'b110;
        rom_memory[7561] = 3'b110;
        rom_memory[7562] = 3'b110;
        rom_memory[7563] = 3'b110;
        rom_memory[7564] = 3'b110;
        rom_memory[7565] = 3'b110;
        rom_memory[7566] = 3'b110;
        rom_memory[7567] = 3'b110;
        rom_memory[7568] = 3'b110;
        rom_memory[7569] = 3'b110;
        rom_memory[7570] = 3'b110;
        rom_memory[7571] = 3'b110;
        rom_memory[7572] = 3'b110;
        rom_memory[7573] = 3'b110;
        rom_memory[7574] = 3'b110;
        rom_memory[7575] = 3'b110;
        rom_memory[7576] = 3'b110;
        rom_memory[7577] = 3'b110;
        rom_memory[7578] = 3'b110;
        rom_memory[7579] = 3'b110;
        rom_memory[7580] = 3'b110;
        rom_memory[7581] = 3'b110;
        rom_memory[7582] = 3'b110;
        rom_memory[7583] = 3'b110;
        rom_memory[7584] = 3'b110;
        rom_memory[7585] = 3'b110;
        rom_memory[7586] = 3'b110;
        rom_memory[7587] = 3'b110;
        rom_memory[7588] = 3'b110;
        rom_memory[7589] = 3'b110;
        rom_memory[7590] = 3'b110;
        rom_memory[7591] = 3'b110;
        rom_memory[7592] = 3'b110;
        rom_memory[7593] = 3'b110;
        rom_memory[7594] = 3'b110;
        rom_memory[7595] = 3'b110;
        rom_memory[7596] = 3'b110;
        rom_memory[7597] = 3'b110;
        rom_memory[7598] = 3'b110;
        rom_memory[7599] = 3'b110;
        rom_memory[7600] = 3'b110;
        rom_memory[7601] = 3'b110;
        rom_memory[7602] = 3'b110;
        rom_memory[7603] = 3'b110;
        rom_memory[7604] = 3'b110;
        rom_memory[7605] = 3'b110;
        rom_memory[7606] = 3'b110;
        rom_memory[7607] = 3'b110;
        rom_memory[7608] = 3'b110;
        rom_memory[7609] = 3'b110;
        rom_memory[7610] = 3'b110;
        rom_memory[7611] = 3'b110;
        rom_memory[7612] = 3'b110;
        rom_memory[7613] = 3'b110;
        rom_memory[7614] = 3'b110;
        rom_memory[7615] = 3'b110;
        rom_memory[7616] = 3'b110;
        rom_memory[7617] = 3'b110;
        rom_memory[7618] = 3'b110;
        rom_memory[7619] = 3'b110;
        rom_memory[7620] = 3'b110;
        rom_memory[7621] = 3'b110;
        rom_memory[7622] = 3'b110;
        rom_memory[7623] = 3'b110;
        rom_memory[7624] = 3'b110;
        rom_memory[7625] = 3'b110;
        rom_memory[7626] = 3'b110;
        rom_memory[7627] = 3'b110;
        rom_memory[7628] = 3'b110;
        rom_memory[7629] = 3'b110;
        rom_memory[7630] = 3'b110;
        rom_memory[7631] = 3'b110;
        rom_memory[7632] = 3'b110;
        rom_memory[7633] = 3'b110;
        rom_memory[7634] = 3'b110;
        rom_memory[7635] = 3'b110;
        rom_memory[7636] = 3'b110;
        rom_memory[7637] = 3'b110;
        rom_memory[7638] = 3'b110;
        rom_memory[7639] = 3'b110;
        rom_memory[7640] = 3'b110;
        rom_memory[7641] = 3'b110;
        rom_memory[7642] = 3'b110;
        rom_memory[7643] = 3'b110;
        rom_memory[7644] = 3'b110;
        rom_memory[7645] = 3'b110;
        rom_memory[7646] = 3'b110;
        rom_memory[7647] = 3'b110;
        rom_memory[7648] = 3'b110;
        rom_memory[7649] = 3'b110;
        rom_memory[7650] = 3'b110;
        rom_memory[7651] = 3'b110;
        rom_memory[7652] = 3'b110;
        rom_memory[7653] = 3'b110;
        rom_memory[7654] = 3'b110;
        rom_memory[7655] = 3'b110;
        rom_memory[7656] = 3'b110;
        rom_memory[7657] = 3'b110;
        rom_memory[7658] = 3'b110;
        rom_memory[7659] = 3'b110;
        rom_memory[7660] = 3'b110;
        rom_memory[7661] = 3'b110;
        rom_memory[7662] = 3'b110;
        rom_memory[7663] = 3'b110;
        rom_memory[7664] = 3'b110;
        rom_memory[7665] = 3'b110;
        rom_memory[7666] = 3'b110;
        rom_memory[7667] = 3'b110;
        rom_memory[7668] = 3'b110;
        rom_memory[7669] = 3'b110;
        rom_memory[7670] = 3'b110;
        rom_memory[7671] = 3'b110;
        rom_memory[7672] = 3'b110;
        rom_memory[7673] = 3'b110;
        rom_memory[7674] = 3'b110;
        rom_memory[7675] = 3'b110;
        rom_memory[7676] = 3'b110;
        rom_memory[7677] = 3'b110;
        rom_memory[7678] = 3'b110;
        rom_memory[7679] = 3'b110;
        rom_memory[7680] = 3'b110;
        rom_memory[7681] = 3'b110;
        rom_memory[7682] = 3'b110;
        rom_memory[7683] = 3'b110;
        rom_memory[7684] = 3'b110;
        rom_memory[7685] = 3'b110;
        rom_memory[7686] = 3'b110;
        rom_memory[7687] = 3'b110;
        rom_memory[7688] = 3'b110;
        rom_memory[7689] = 3'b110;
        rom_memory[7690] = 3'b110;
        rom_memory[7691] = 3'b110;
        rom_memory[7692] = 3'b110;
        rom_memory[7693] = 3'b110;
        rom_memory[7694] = 3'b110;
        rom_memory[7695] = 3'b110;
        rom_memory[7696] = 3'b110;
        rom_memory[7697] = 3'b110;
        rom_memory[7698] = 3'b110;
        rom_memory[7699] = 3'b110;
        rom_memory[7700] = 3'b110;
        rom_memory[7701] = 3'b110;
        rom_memory[7702] = 3'b110;
        rom_memory[7703] = 3'b110;
        rom_memory[7704] = 3'b110;
        rom_memory[7705] = 3'b110;
        rom_memory[7706] = 3'b110;
        rom_memory[7707] = 3'b110;
        rom_memory[7708] = 3'b110;
        rom_memory[7709] = 3'b110;
        rom_memory[7710] = 3'b110;
        rom_memory[7711] = 3'b110;
        rom_memory[7712] = 3'b110;
        rom_memory[7713] = 3'b110;
        rom_memory[7714] = 3'b110;
        rom_memory[7715] = 3'b110;
        rom_memory[7716] = 3'b110;
        rom_memory[7717] = 3'b110;
        rom_memory[7718] = 3'b110;
        rom_memory[7719] = 3'b110;
        rom_memory[7720] = 3'b110;
        rom_memory[7721] = 3'b110;
        rom_memory[7722] = 3'b110;
        rom_memory[7723] = 3'b110;
        rom_memory[7724] = 3'b110;
        rom_memory[7725] = 3'b000;
        rom_memory[7726] = 3'b000;
        rom_memory[7727] = 3'b000;
        rom_memory[7728] = 3'b100;
        rom_memory[7729] = 3'b111;
        rom_memory[7730] = 3'b111;
        rom_memory[7731] = 3'b111;
        rom_memory[7732] = 3'b000;
        rom_memory[7733] = 3'b000;
        rom_memory[7734] = 3'b000;
        rom_memory[7735] = 3'b000;
        rom_memory[7736] = 3'b000;
        rom_memory[7737] = 3'b000;
        rom_memory[7738] = 3'b000;
        rom_memory[7739] = 3'b000;
        rom_memory[7740] = 3'b000;
        rom_memory[7741] = 3'b000;
        rom_memory[7742] = 3'b000;
        rom_memory[7743] = 3'b000;
        rom_memory[7744] = 3'b000;
        rom_memory[7745] = 3'b000;
        rom_memory[7746] = 3'b000;
        rom_memory[7747] = 3'b000;
        rom_memory[7748] = 3'b000;
        rom_memory[7749] = 3'b000;
        rom_memory[7750] = 3'b000;
        rom_memory[7751] = 3'b000;
        rom_memory[7752] = 3'b000;
        rom_memory[7753] = 3'b000;
        rom_memory[7754] = 3'b000;
        rom_memory[7755] = 3'b000;
        rom_memory[7756] = 3'b011;
        rom_memory[7757] = 3'b011;
        rom_memory[7758] = 3'b000;
        rom_memory[7759] = 3'b000;
        rom_memory[7760] = 3'b000;
        rom_memory[7761] = 3'b010;
        rom_memory[7762] = 3'b010;
        rom_memory[7763] = 3'b000;
        rom_memory[7764] = 3'b011;
        rom_memory[7765] = 3'b011;
        rom_memory[7766] = 3'b011;
        rom_memory[7767] = 3'b001;
        rom_memory[7768] = 3'b001;
        rom_memory[7769] = 3'b001;
        rom_memory[7770] = 3'b111;
        rom_memory[7771] = 3'b111;
        rom_memory[7772] = 3'b111;
        rom_memory[7773] = 3'b110;
        rom_memory[7774] = 3'b110;
        rom_memory[7775] = 3'b110;
        rom_memory[7776] = 3'b110;
        rom_memory[7777] = 3'b110;
        rom_memory[7778] = 3'b110;
        rom_memory[7779] = 3'b110;
        rom_memory[7780] = 3'b110;
        rom_memory[7781] = 3'b110;
        rom_memory[7782] = 3'b110;
        rom_memory[7783] = 3'b110;
        rom_memory[7784] = 3'b110;
        rom_memory[7785] = 3'b110;
        rom_memory[7786] = 3'b110;
        rom_memory[7787] = 3'b110;
        rom_memory[7788] = 3'b110;
        rom_memory[7789] = 3'b110;
        rom_memory[7790] = 3'b110;
        rom_memory[7791] = 3'b110;
        rom_memory[7792] = 3'b110;
        rom_memory[7793] = 3'b110;
        rom_memory[7794] = 3'b110;
        rom_memory[7795] = 3'b110;
        rom_memory[7796] = 3'b110;
        rom_memory[7797] = 3'b110;
        rom_memory[7798] = 3'b110;
        rom_memory[7799] = 3'b110;
        rom_memory[7800] = 3'b110;
        rom_memory[7801] = 3'b110;
        rom_memory[7802] = 3'b110;
        rom_memory[7803] = 3'b110;
        rom_memory[7804] = 3'b110;
        rom_memory[7805] = 3'b110;
        rom_memory[7806] = 3'b110;
        rom_memory[7807] = 3'b110;
        rom_memory[7808] = 3'b110;
        rom_memory[7809] = 3'b110;
        rom_memory[7810] = 3'b110;
        rom_memory[7811] = 3'b110;
        rom_memory[7812] = 3'b110;
        rom_memory[7813] = 3'b110;
        rom_memory[7814] = 3'b110;
        rom_memory[7815] = 3'b110;
        rom_memory[7816] = 3'b110;
        rom_memory[7817] = 3'b110;
        rom_memory[7818] = 3'b110;
        rom_memory[7819] = 3'b110;
        rom_memory[7820] = 3'b110;
        rom_memory[7821] = 3'b110;
        rom_memory[7822] = 3'b110;
        rom_memory[7823] = 3'b110;
        rom_memory[7824] = 3'b110;
        rom_memory[7825] = 3'b110;
        rom_memory[7826] = 3'b110;
        rom_memory[7827] = 3'b110;
        rom_memory[7828] = 3'b110;
        rom_memory[7829] = 3'b110;
        rom_memory[7830] = 3'b110;
        rom_memory[7831] = 3'b110;
        rom_memory[7832] = 3'b110;
        rom_memory[7833] = 3'b110;
        rom_memory[7834] = 3'b110;
        rom_memory[7835] = 3'b110;
        rom_memory[7836] = 3'b110;
        rom_memory[7837] = 3'b110;
        rom_memory[7838] = 3'b110;
        rom_memory[7839] = 3'b110;
        rom_memory[7840] = 3'b110;
        rom_memory[7841] = 3'b110;
        rom_memory[7842] = 3'b110;
        rom_memory[7843] = 3'b110;
        rom_memory[7844] = 3'b110;
        rom_memory[7845] = 3'b110;
        rom_memory[7846] = 3'b110;
        rom_memory[7847] = 3'b110;
        rom_memory[7848] = 3'b110;
        rom_memory[7849] = 3'b110;
        rom_memory[7850] = 3'b110;
        rom_memory[7851] = 3'b110;
        rom_memory[7852] = 3'b110;
        rom_memory[7853] = 3'b110;
        rom_memory[7854] = 3'b110;
        rom_memory[7855] = 3'b110;
        rom_memory[7856] = 3'b110;
        rom_memory[7857] = 3'b110;
        rom_memory[7858] = 3'b110;
        rom_memory[7859] = 3'b110;
        rom_memory[7860] = 3'b110;
        rom_memory[7861] = 3'b110;
        rom_memory[7862] = 3'b110;
        rom_memory[7863] = 3'b110;
        rom_memory[7864] = 3'b110;
        rom_memory[7865] = 3'b110;
        rom_memory[7866] = 3'b110;
        rom_memory[7867] = 3'b110;
        rom_memory[7868] = 3'b110;
        rom_memory[7869] = 3'b110;
        rom_memory[7870] = 3'b110;
        rom_memory[7871] = 3'b110;
        rom_memory[7872] = 3'b110;
        rom_memory[7873] = 3'b110;
        rom_memory[7874] = 3'b110;
        rom_memory[7875] = 3'b110;
        rom_memory[7876] = 3'b110;
        rom_memory[7877] = 3'b110;
        rom_memory[7878] = 3'b110;
        rom_memory[7879] = 3'b110;
        rom_memory[7880] = 3'b110;
        rom_memory[7881] = 3'b110;
        rom_memory[7882] = 3'b110;
        rom_memory[7883] = 3'b110;
        rom_memory[7884] = 3'b110;
        rom_memory[7885] = 3'b110;
        rom_memory[7886] = 3'b110;
        rom_memory[7887] = 3'b110;
        rom_memory[7888] = 3'b110;
        rom_memory[7889] = 3'b110;
        rom_memory[7890] = 3'b110;
        rom_memory[7891] = 3'b110;
        rom_memory[7892] = 3'b110;
        rom_memory[7893] = 3'b110;
        rom_memory[7894] = 3'b110;
        rom_memory[7895] = 3'b110;
        rom_memory[7896] = 3'b110;
        rom_memory[7897] = 3'b110;
        rom_memory[7898] = 3'b110;
        rom_memory[7899] = 3'b110;
        rom_memory[7900] = 3'b110;
        rom_memory[7901] = 3'b110;
        rom_memory[7902] = 3'b110;
        rom_memory[7903] = 3'b110;
        rom_memory[7904] = 3'b110;
        rom_memory[7905] = 3'b110;
        rom_memory[7906] = 3'b110;
        rom_memory[7907] = 3'b110;
        rom_memory[7908] = 3'b110;
        rom_memory[7909] = 3'b110;
        rom_memory[7910] = 3'b110;
        rom_memory[7911] = 3'b110;
        rom_memory[7912] = 3'b110;
        rom_memory[7913] = 3'b110;
        rom_memory[7914] = 3'b110;
        rom_memory[7915] = 3'b110;
        rom_memory[7916] = 3'b110;
        rom_memory[7917] = 3'b110;
        rom_memory[7918] = 3'b110;
        rom_memory[7919] = 3'b110;
        rom_memory[7920] = 3'b110;
        rom_memory[7921] = 3'b110;
        rom_memory[7922] = 3'b110;
        rom_memory[7923] = 3'b110;
        rom_memory[7924] = 3'b110;
        rom_memory[7925] = 3'b110;
        rom_memory[7926] = 3'b110;
        rom_memory[7927] = 3'b110;
        rom_memory[7928] = 3'b110;
        rom_memory[7929] = 3'b110;
        rom_memory[7930] = 3'b110;
        rom_memory[7931] = 3'b110;
        rom_memory[7932] = 3'b110;
        rom_memory[7933] = 3'b110;
        rom_memory[7934] = 3'b110;
        rom_memory[7935] = 3'b110;
        rom_memory[7936] = 3'b110;
        rom_memory[7937] = 3'b110;
        rom_memory[7938] = 3'b110;
        rom_memory[7939] = 3'b110;
        rom_memory[7940] = 3'b110;
        rom_memory[7941] = 3'b110;
        rom_memory[7942] = 3'b110;
        rom_memory[7943] = 3'b110;
        rom_memory[7944] = 3'b110;
        rom_memory[7945] = 3'b110;
        rom_memory[7946] = 3'b110;
        rom_memory[7947] = 3'b110;
        rom_memory[7948] = 3'b110;
        rom_memory[7949] = 3'b110;
        rom_memory[7950] = 3'b110;
        rom_memory[7951] = 3'b110;
        rom_memory[7952] = 3'b110;
        rom_memory[7953] = 3'b110;
        rom_memory[7954] = 3'b110;
        rom_memory[7955] = 3'b110;
        rom_memory[7956] = 3'b110;
        rom_memory[7957] = 3'b110;
        rom_memory[7958] = 3'b110;
        rom_memory[7959] = 3'b110;
        rom_memory[7960] = 3'b110;
        rom_memory[7961] = 3'b110;
        rom_memory[7962] = 3'b110;
        rom_memory[7963] = 3'b110;
        rom_memory[7964] = 3'b110;
        rom_memory[7965] = 3'b000;
        rom_memory[7966] = 3'b000;
        rom_memory[7967] = 3'b000;
        rom_memory[7968] = 3'b000;
        rom_memory[7969] = 3'b100;
        rom_memory[7970] = 3'b100;
        rom_memory[7971] = 3'b111;
        rom_memory[7972] = 3'b111;
        rom_memory[7973] = 3'b000;
        rom_memory[7974] = 3'b000;
        rom_memory[7975] = 3'b000;
        rom_memory[7976] = 3'b000;
        rom_memory[7977] = 3'b000;
        rom_memory[7978] = 3'b000;
        rom_memory[7979] = 3'b000;
        rom_memory[7980] = 3'b000;
        rom_memory[7981] = 3'b000;
        rom_memory[7982] = 3'b000;
        rom_memory[7983] = 3'b000;
        rom_memory[7984] = 3'b000;
        rom_memory[7985] = 3'b000;
        rom_memory[7986] = 3'b000;
        rom_memory[7987] = 3'b000;
        rom_memory[7988] = 3'b000;
        rom_memory[7989] = 3'b000;
        rom_memory[7990] = 3'b000;
        rom_memory[7991] = 3'b000;
        rom_memory[7992] = 3'b000;
        rom_memory[7993] = 3'b000;
        rom_memory[7994] = 3'b000;
        rom_memory[7995] = 3'b000;
        rom_memory[7996] = 3'b000;
        rom_memory[7997] = 3'b000;
        rom_memory[7998] = 3'b000;
        rom_memory[7999] = 3'b010;
        rom_memory[8000] = 3'b010;
        rom_memory[8001] = 3'b010;
        rom_memory[8002] = 3'b011;
        rom_memory[8003] = 3'b011;
        rom_memory[8004] = 3'b011;
        rom_memory[8005] = 3'b011;
        rom_memory[8006] = 3'b011;
        rom_memory[8007] = 3'b011;
        rom_memory[8008] = 3'b011;
        rom_memory[8009] = 3'b011;
        rom_memory[8010] = 3'b011;
        rom_memory[8011] = 3'b111;
        rom_memory[8012] = 3'b111;
        rom_memory[8013] = 3'b111;
        rom_memory[8014] = 3'b110;
        rom_memory[8015] = 3'b110;
        rom_memory[8016] = 3'b110;
        rom_memory[8017] = 3'b110;
        rom_memory[8018] = 3'b110;
        rom_memory[8019] = 3'b110;
        rom_memory[8020] = 3'b110;
        rom_memory[8021] = 3'b110;
        rom_memory[8022] = 3'b110;
        rom_memory[8023] = 3'b110;
        rom_memory[8024] = 3'b110;
        rom_memory[8025] = 3'b110;
        rom_memory[8026] = 3'b110;
        rom_memory[8027] = 3'b110;
        rom_memory[8028] = 3'b110;
        rom_memory[8029] = 3'b110;
        rom_memory[8030] = 3'b110;
        rom_memory[8031] = 3'b110;
        rom_memory[8032] = 3'b110;
        rom_memory[8033] = 3'b110;
        rom_memory[8034] = 3'b110;
        rom_memory[8035] = 3'b110;
        rom_memory[8036] = 3'b110;
        rom_memory[8037] = 3'b110;
        rom_memory[8038] = 3'b110;
        rom_memory[8039] = 3'b110;
        rom_memory[8040] = 3'b110;
        rom_memory[8041] = 3'b110;
        rom_memory[8042] = 3'b110;
        rom_memory[8043] = 3'b110;
        rom_memory[8044] = 3'b110;
        rom_memory[8045] = 3'b110;
        rom_memory[8046] = 3'b110;
        rom_memory[8047] = 3'b110;
        rom_memory[8048] = 3'b110;
        rom_memory[8049] = 3'b110;
        rom_memory[8050] = 3'b110;
        rom_memory[8051] = 3'b110;
        rom_memory[8052] = 3'b110;
        rom_memory[8053] = 3'b110;
        rom_memory[8054] = 3'b110;
        rom_memory[8055] = 3'b110;
        rom_memory[8056] = 3'b110;
        rom_memory[8057] = 3'b110;
        rom_memory[8058] = 3'b110;
        rom_memory[8059] = 3'b110;
        rom_memory[8060] = 3'b110;
        rom_memory[8061] = 3'b110;
        rom_memory[8062] = 3'b110;
        rom_memory[8063] = 3'b110;
        rom_memory[8064] = 3'b110;
        rom_memory[8065] = 3'b110;
        rom_memory[8066] = 3'b110;
        rom_memory[8067] = 3'b110;
        rom_memory[8068] = 3'b110;
        rom_memory[8069] = 3'b110;
        rom_memory[8070] = 3'b110;
        rom_memory[8071] = 3'b110;
        rom_memory[8072] = 3'b110;
        rom_memory[8073] = 3'b110;
        rom_memory[8074] = 3'b110;
        rom_memory[8075] = 3'b110;
        rom_memory[8076] = 3'b110;
        rom_memory[8077] = 3'b110;
        rom_memory[8078] = 3'b110;
        rom_memory[8079] = 3'b110;
        rom_memory[8080] = 3'b110;
        rom_memory[8081] = 3'b110;
        rom_memory[8082] = 3'b110;
        rom_memory[8083] = 3'b110;
        rom_memory[8084] = 3'b110;
        rom_memory[8085] = 3'b110;
        rom_memory[8086] = 3'b110;
        rom_memory[8087] = 3'b110;
        rom_memory[8088] = 3'b110;
        rom_memory[8089] = 3'b110;
        rom_memory[8090] = 3'b110;
        rom_memory[8091] = 3'b110;
        rom_memory[8092] = 3'b110;
        rom_memory[8093] = 3'b110;
        rom_memory[8094] = 3'b110;
        rom_memory[8095] = 3'b110;
        rom_memory[8096] = 3'b110;
        rom_memory[8097] = 3'b110;
        rom_memory[8098] = 3'b110;
        rom_memory[8099] = 3'b110;
        rom_memory[8100] = 3'b110;
        rom_memory[8101] = 3'b110;
        rom_memory[8102] = 3'b110;
        rom_memory[8103] = 3'b110;
        rom_memory[8104] = 3'b110;
        rom_memory[8105] = 3'b110;
        rom_memory[8106] = 3'b110;
        rom_memory[8107] = 3'b110;
        rom_memory[8108] = 3'b110;
        rom_memory[8109] = 3'b110;
        rom_memory[8110] = 3'b110;
        rom_memory[8111] = 3'b110;
        rom_memory[8112] = 3'b110;
        rom_memory[8113] = 3'b110;
        rom_memory[8114] = 3'b110;
        rom_memory[8115] = 3'b110;
        rom_memory[8116] = 3'b110;
        rom_memory[8117] = 3'b110;
        rom_memory[8118] = 3'b110;
        rom_memory[8119] = 3'b110;
        rom_memory[8120] = 3'b110;
        rom_memory[8121] = 3'b110;
        rom_memory[8122] = 3'b110;
        rom_memory[8123] = 3'b110;
        rom_memory[8124] = 3'b110;
        rom_memory[8125] = 3'b110;
        rom_memory[8126] = 3'b110;
        rom_memory[8127] = 3'b110;
        rom_memory[8128] = 3'b110;
        rom_memory[8129] = 3'b110;
        rom_memory[8130] = 3'b110;
        rom_memory[8131] = 3'b110;
        rom_memory[8132] = 3'b110;
        rom_memory[8133] = 3'b110;
        rom_memory[8134] = 3'b110;
        rom_memory[8135] = 3'b110;
        rom_memory[8136] = 3'b110;
        rom_memory[8137] = 3'b110;
        rom_memory[8138] = 3'b110;
        rom_memory[8139] = 3'b110;
        rom_memory[8140] = 3'b110;
        rom_memory[8141] = 3'b110;
        rom_memory[8142] = 3'b110;
        rom_memory[8143] = 3'b110;
        rom_memory[8144] = 3'b110;
        rom_memory[8145] = 3'b110;
        rom_memory[8146] = 3'b110;
        rom_memory[8147] = 3'b110;
        rom_memory[8148] = 3'b110;
        rom_memory[8149] = 3'b110;
        rom_memory[8150] = 3'b110;
        rom_memory[8151] = 3'b110;
        rom_memory[8152] = 3'b110;
        rom_memory[8153] = 3'b110;
        rom_memory[8154] = 3'b110;
        rom_memory[8155] = 3'b110;
        rom_memory[8156] = 3'b110;
        rom_memory[8157] = 3'b110;
        rom_memory[8158] = 3'b110;
        rom_memory[8159] = 3'b110;
        rom_memory[8160] = 3'b110;
        rom_memory[8161] = 3'b110;
        rom_memory[8162] = 3'b110;
        rom_memory[8163] = 3'b110;
        rom_memory[8164] = 3'b110;
        rom_memory[8165] = 3'b110;
        rom_memory[8166] = 3'b110;
        rom_memory[8167] = 3'b110;
        rom_memory[8168] = 3'b110;
        rom_memory[8169] = 3'b110;
        rom_memory[8170] = 3'b110;
        rom_memory[8171] = 3'b110;
        rom_memory[8172] = 3'b110;
        rom_memory[8173] = 3'b110;
        rom_memory[8174] = 3'b110;
        rom_memory[8175] = 3'b110;
        rom_memory[8176] = 3'b110;
        rom_memory[8177] = 3'b110;
        rom_memory[8178] = 3'b110;
        rom_memory[8179] = 3'b110;
        rom_memory[8180] = 3'b110;
        rom_memory[8181] = 3'b110;
        rom_memory[8182] = 3'b110;
        rom_memory[8183] = 3'b110;
        rom_memory[8184] = 3'b110;
        rom_memory[8185] = 3'b110;
        rom_memory[8186] = 3'b110;
        rom_memory[8187] = 3'b110;
        rom_memory[8188] = 3'b110;
        rom_memory[8189] = 3'b110;
        rom_memory[8190] = 3'b110;
        rom_memory[8191] = 3'b110;
        rom_memory[8192] = 3'b110;
        rom_memory[8193] = 3'b110;
        rom_memory[8194] = 3'b110;
        rom_memory[8195] = 3'b110;
        rom_memory[8196] = 3'b110;
        rom_memory[8197] = 3'b110;
        rom_memory[8198] = 3'b110;
        rom_memory[8199] = 3'b110;
        rom_memory[8200] = 3'b110;
        rom_memory[8201] = 3'b110;
        rom_memory[8202] = 3'b110;
        rom_memory[8203] = 3'b110;
        rom_memory[8204] = 3'b110;
        rom_memory[8205] = 3'b100;
        rom_memory[8206] = 3'b000;
        rom_memory[8207] = 3'b000;
        rom_memory[8208] = 3'b000;
        rom_memory[8209] = 3'b000;
        rom_memory[8210] = 3'b000;
        rom_memory[8211] = 3'b000;
        rom_memory[8212] = 3'b000;
        rom_memory[8213] = 3'b000;
        rom_memory[8214] = 3'b000;
        rom_memory[8215] = 3'b000;
        rom_memory[8216] = 3'b000;
        rom_memory[8217] = 3'b000;
        rom_memory[8218] = 3'b000;
        rom_memory[8219] = 3'b000;
        rom_memory[8220] = 3'b000;
        rom_memory[8221] = 3'b000;
        rom_memory[8222] = 3'b000;
        rom_memory[8223] = 3'b000;
        rom_memory[8224] = 3'b000;
        rom_memory[8225] = 3'b000;
        rom_memory[8226] = 3'b000;
        rom_memory[8227] = 3'b000;
        rom_memory[8228] = 3'b000;
        rom_memory[8229] = 3'b000;
        rom_memory[8230] = 3'b000;
        rom_memory[8231] = 3'b000;
        rom_memory[8232] = 3'b000;
        rom_memory[8233] = 3'b000;
        rom_memory[8234] = 3'b000;
        rom_memory[8235] = 3'b000;
        rom_memory[8236] = 3'b000;
        rom_memory[8237] = 3'b000;
        rom_memory[8238] = 3'b010;
        rom_memory[8239] = 3'b010;
        rom_memory[8240] = 3'b010;
        rom_memory[8241] = 3'b010;
        rom_memory[8242] = 3'b010;
        rom_memory[8243] = 3'b011;
        rom_memory[8244] = 3'b011;
        rom_memory[8245] = 3'b011;
        rom_memory[8246] = 3'b011;
        rom_memory[8247] = 3'b011;
        rom_memory[8248] = 3'b011;
        rom_memory[8249] = 3'b011;
        rom_memory[8250] = 3'b001;
        rom_memory[8251] = 3'b011;
        rom_memory[8252] = 3'b111;
        rom_memory[8253] = 3'b111;
        rom_memory[8254] = 3'b110;
        rom_memory[8255] = 3'b110;
        rom_memory[8256] = 3'b110;
        rom_memory[8257] = 3'b110;
        rom_memory[8258] = 3'b110;
        rom_memory[8259] = 3'b110;
        rom_memory[8260] = 3'b110;
        rom_memory[8261] = 3'b110;
        rom_memory[8262] = 3'b110;
        rom_memory[8263] = 3'b110;
        rom_memory[8264] = 3'b110;
        rom_memory[8265] = 3'b110;
        rom_memory[8266] = 3'b110;
        rom_memory[8267] = 3'b110;
        rom_memory[8268] = 3'b110;
        rom_memory[8269] = 3'b110;
        rom_memory[8270] = 3'b110;
        rom_memory[8271] = 3'b110;
        rom_memory[8272] = 3'b110;
        rom_memory[8273] = 3'b110;
        rom_memory[8274] = 3'b110;
        rom_memory[8275] = 3'b110;
        rom_memory[8276] = 3'b110;
        rom_memory[8277] = 3'b110;
        rom_memory[8278] = 3'b110;
        rom_memory[8279] = 3'b110;
        rom_memory[8280] = 3'b110;
        rom_memory[8281] = 3'b110;
        rom_memory[8282] = 3'b110;
        rom_memory[8283] = 3'b110;
        rom_memory[8284] = 3'b110;
        rom_memory[8285] = 3'b110;
        rom_memory[8286] = 3'b110;
        rom_memory[8287] = 3'b110;
        rom_memory[8288] = 3'b110;
        rom_memory[8289] = 3'b110;
        rom_memory[8290] = 3'b110;
        rom_memory[8291] = 3'b110;
        rom_memory[8292] = 3'b110;
        rom_memory[8293] = 3'b110;
        rom_memory[8294] = 3'b110;
        rom_memory[8295] = 3'b110;
        rom_memory[8296] = 3'b110;
        rom_memory[8297] = 3'b110;
        rom_memory[8298] = 3'b110;
        rom_memory[8299] = 3'b110;
        rom_memory[8300] = 3'b110;
        rom_memory[8301] = 3'b110;
        rom_memory[8302] = 3'b110;
        rom_memory[8303] = 3'b110;
        rom_memory[8304] = 3'b110;
        rom_memory[8305] = 3'b110;
        rom_memory[8306] = 3'b110;
        rom_memory[8307] = 3'b110;
        rom_memory[8308] = 3'b110;
        rom_memory[8309] = 3'b110;
        rom_memory[8310] = 3'b110;
        rom_memory[8311] = 3'b110;
        rom_memory[8312] = 3'b110;
        rom_memory[8313] = 3'b110;
        rom_memory[8314] = 3'b110;
        rom_memory[8315] = 3'b110;
        rom_memory[8316] = 3'b110;
        rom_memory[8317] = 3'b110;
        rom_memory[8318] = 3'b110;
        rom_memory[8319] = 3'b110;
        rom_memory[8320] = 3'b110;
        rom_memory[8321] = 3'b110;
        rom_memory[8322] = 3'b110;
        rom_memory[8323] = 3'b110;
        rom_memory[8324] = 3'b110;
        rom_memory[8325] = 3'b110;
        rom_memory[8326] = 3'b110;
        rom_memory[8327] = 3'b110;
        rom_memory[8328] = 3'b110;
        rom_memory[8329] = 3'b110;
        rom_memory[8330] = 3'b110;
        rom_memory[8331] = 3'b110;
        rom_memory[8332] = 3'b110;
        rom_memory[8333] = 3'b110;
        rom_memory[8334] = 3'b110;
        rom_memory[8335] = 3'b110;
        rom_memory[8336] = 3'b110;
        rom_memory[8337] = 3'b110;
        rom_memory[8338] = 3'b110;
        rom_memory[8339] = 3'b110;
        rom_memory[8340] = 3'b110;
        rom_memory[8341] = 3'b110;
        rom_memory[8342] = 3'b110;
        rom_memory[8343] = 3'b110;
        rom_memory[8344] = 3'b110;
        rom_memory[8345] = 3'b110;
        rom_memory[8346] = 3'b110;
        rom_memory[8347] = 3'b110;
        rom_memory[8348] = 3'b110;
        rom_memory[8349] = 3'b110;
        rom_memory[8350] = 3'b110;
        rom_memory[8351] = 3'b110;
        rom_memory[8352] = 3'b110;
        rom_memory[8353] = 3'b110;
        rom_memory[8354] = 3'b110;
        rom_memory[8355] = 3'b110;
        rom_memory[8356] = 3'b110;
        rom_memory[8357] = 3'b110;
        rom_memory[8358] = 3'b110;
        rom_memory[8359] = 3'b110;
        rom_memory[8360] = 3'b110;
        rom_memory[8361] = 3'b110;
        rom_memory[8362] = 3'b110;
        rom_memory[8363] = 3'b110;
        rom_memory[8364] = 3'b110;
        rom_memory[8365] = 3'b110;
        rom_memory[8366] = 3'b110;
        rom_memory[8367] = 3'b110;
        rom_memory[8368] = 3'b110;
        rom_memory[8369] = 3'b110;
        rom_memory[8370] = 3'b110;
        rom_memory[8371] = 3'b110;
        rom_memory[8372] = 3'b110;
        rom_memory[8373] = 3'b110;
        rom_memory[8374] = 3'b110;
        rom_memory[8375] = 3'b110;
        rom_memory[8376] = 3'b110;
        rom_memory[8377] = 3'b110;
        rom_memory[8378] = 3'b110;
        rom_memory[8379] = 3'b110;
        rom_memory[8380] = 3'b110;
        rom_memory[8381] = 3'b110;
        rom_memory[8382] = 3'b110;
        rom_memory[8383] = 3'b110;
        rom_memory[8384] = 3'b110;
        rom_memory[8385] = 3'b110;
        rom_memory[8386] = 3'b110;
        rom_memory[8387] = 3'b110;
        rom_memory[8388] = 3'b110;
        rom_memory[8389] = 3'b110;
        rom_memory[8390] = 3'b110;
        rom_memory[8391] = 3'b110;
        rom_memory[8392] = 3'b110;
        rom_memory[8393] = 3'b110;
        rom_memory[8394] = 3'b110;
        rom_memory[8395] = 3'b110;
        rom_memory[8396] = 3'b110;
        rom_memory[8397] = 3'b110;
        rom_memory[8398] = 3'b110;
        rom_memory[8399] = 3'b110;
        rom_memory[8400] = 3'b110;
        rom_memory[8401] = 3'b110;
        rom_memory[8402] = 3'b110;
        rom_memory[8403] = 3'b110;
        rom_memory[8404] = 3'b110;
        rom_memory[8405] = 3'b110;
        rom_memory[8406] = 3'b110;
        rom_memory[8407] = 3'b110;
        rom_memory[8408] = 3'b110;
        rom_memory[8409] = 3'b110;
        rom_memory[8410] = 3'b110;
        rom_memory[8411] = 3'b110;
        rom_memory[8412] = 3'b110;
        rom_memory[8413] = 3'b110;
        rom_memory[8414] = 3'b110;
        rom_memory[8415] = 3'b110;
        rom_memory[8416] = 3'b110;
        rom_memory[8417] = 3'b110;
        rom_memory[8418] = 3'b110;
        rom_memory[8419] = 3'b110;
        rom_memory[8420] = 3'b110;
        rom_memory[8421] = 3'b110;
        rom_memory[8422] = 3'b110;
        rom_memory[8423] = 3'b110;
        rom_memory[8424] = 3'b110;
        rom_memory[8425] = 3'b110;
        rom_memory[8426] = 3'b110;
        rom_memory[8427] = 3'b110;
        rom_memory[8428] = 3'b110;
        rom_memory[8429] = 3'b110;
        rom_memory[8430] = 3'b110;
        rom_memory[8431] = 3'b110;
        rom_memory[8432] = 3'b110;
        rom_memory[8433] = 3'b110;
        rom_memory[8434] = 3'b110;
        rom_memory[8435] = 3'b110;
        rom_memory[8436] = 3'b110;
        rom_memory[8437] = 3'b110;
        rom_memory[8438] = 3'b110;
        rom_memory[8439] = 3'b110;
        rom_memory[8440] = 3'b110;
        rom_memory[8441] = 3'b110;
        rom_memory[8442] = 3'b110;
        rom_memory[8443] = 3'b110;
        rom_memory[8444] = 3'b110;
        rom_memory[8445] = 3'b110;
        rom_memory[8446] = 3'b000;
        rom_memory[8447] = 3'b000;
        rom_memory[8448] = 3'b000;
        rom_memory[8449] = 3'b000;
        rom_memory[8450] = 3'b000;
        rom_memory[8451] = 3'b000;
        rom_memory[8452] = 3'b000;
        rom_memory[8453] = 3'b000;
        rom_memory[8454] = 3'b000;
        rom_memory[8455] = 3'b000;
        rom_memory[8456] = 3'b000;
        rom_memory[8457] = 3'b000;
        rom_memory[8458] = 3'b000;
        rom_memory[8459] = 3'b000;
        rom_memory[8460] = 3'b000;
        rom_memory[8461] = 3'b000;
        rom_memory[8462] = 3'b000;
        rom_memory[8463] = 3'b001;
        rom_memory[8464] = 3'b111;
        rom_memory[8465] = 3'b000;
        rom_memory[8466] = 3'b000;
        rom_memory[8467] = 3'b000;
        rom_memory[8468] = 3'b000;
        rom_memory[8469] = 3'b000;
        rom_memory[8470] = 3'b000;
        rom_memory[8471] = 3'b000;
        rom_memory[8472] = 3'b000;
        rom_memory[8473] = 3'b000;
        rom_memory[8474] = 3'b000;
        rom_memory[8475] = 3'b000;
        rom_memory[8476] = 3'b000;
        rom_memory[8477] = 3'b000;
        rom_memory[8478] = 3'b000;
        rom_memory[8479] = 3'b000;
        rom_memory[8480] = 3'b000;
        rom_memory[8481] = 3'b010;
        rom_memory[8482] = 3'b000;
        rom_memory[8483] = 3'b011;
        rom_memory[8484] = 3'b011;
        rom_memory[8485] = 3'b010;
        rom_memory[8486] = 3'b011;
        rom_memory[8487] = 3'b011;
        rom_memory[8488] = 3'b011;
        rom_memory[8489] = 3'b011;
        rom_memory[8490] = 3'b011;
        rom_memory[8491] = 3'b011;
        rom_memory[8492] = 3'b011;
        rom_memory[8493] = 3'b111;
        rom_memory[8494] = 3'b111;
        rom_memory[8495] = 3'b110;
        rom_memory[8496] = 3'b110;
        rom_memory[8497] = 3'b110;
        rom_memory[8498] = 3'b110;
        rom_memory[8499] = 3'b110;
        rom_memory[8500] = 3'b110;
        rom_memory[8501] = 3'b110;
        rom_memory[8502] = 3'b110;
        rom_memory[8503] = 3'b110;
        rom_memory[8504] = 3'b110;
        rom_memory[8505] = 3'b110;
        rom_memory[8506] = 3'b110;
        rom_memory[8507] = 3'b110;
        rom_memory[8508] = 3'b110;
        rom_memory[8509] = 3'b110;
        rom_memory[8510] = 3'b110;
        rom_memory[8511] = 3'b110;
        rom_memory[8512] = 3'b110;
        rom_memory[8513] = 3'b110;
        rom_memory[8514] = 3'b110;
        rom_memory[8515] = 3'b110;
        rom_memory[8516] = 3'b110;
        rom_memory[8517] = 3'b110;
        rom_memory[8518] = 3'b110;
        rom_memory[8519] = 3'b110;
        rom_memory[8520] = 3'b110;
        rom_memory[8521] = 3'b110;
        rom_memory[8522] = 3'b110;
        rom_memory[8523] = 3'b110;
        rom_memory[8524] = 3'b110;
        rom_memory[8525] = 3'b110;
        rom_memory[8526] = 3'b110;
        rom_memory[8527] = 3'b110;
        rom_memory[8528] = 3'b110;
        rom_memory[8529] = 3'b110;
        rom_memory[8530] = 3'b110;
        rom_memory[8531] = 3'b110;
        rom_memory[8532] = 3'b110;
        rom_memory[8533] = 3'b110;
        rom_memory[8534] = 3'b110;
        rom_memory[8535] = 3'b110;
        rom_memory[8536] = 3'b110;
        rom_memory[8537] = 3'b110;
        rom_memory[8538] = 3'b110;
        rom_memory[8539] = 3'b110;
        rom_memory[8540] = 3'b110;
        rom_memory[8541] = 3'b110;
        rom_memory[8542] = 3'b110;
        rom_memory[8543] = 3'b110;
        rom_memory[8544] = 3'b110;
        rom_memory[8545] = 3'b110;
        rom_memory[8546] = 3'b110;
        rom_memory[8547] = 3'b110;
        rom_memory[8548] = 3'b110;
        rom_memory[8549] = 3'b110;
        rom_memory[8550] = 3'b110;
        rom_memory[8551] = 3'b110;
        rom_memory[8552] = 3'b110;
        rom_memory[8553] = 3'b110;
        rom_memory[8554] = 3'b110;
        rom_memory[8555] = 3'b110;
        rom_memory[8556] = 3'b110;
        rom_memory[8557] = 3'b110;
        rom_memory[8558] = 3'b110;
        rom_memory[8559] = 3'b110;
        rom_memory[8560] = 3'b110;
        rom_memory[8561] = 3'b110;
        rom_memory[8562] = 3'b110;
        rom_memory[8563] = 3'b110;
        rom_memory[8564] = 3'b110;
        rom_memory[8565] = 3'b110;
        rom_memory[8566] = 3'b110;
        rom_memory[8567] = 3'b110;
        rom_memory[8568] = 3'b110;
        rom_memory[8569] = 3'b110;
        rom_memory[8570] = 3'b110;
        rom_memory[8571] = 3'b110;
        rom_memory[8572] = 3'b110;
        rom_memory[8573] = 3'b110;
        rom_memory[8574] = 3'b110;
        rom_memory[8575] = 3'b110;
        rom_memory[8576] = 3'b110;
        rom_memory[8577] = 3'b110;
        rom_memory[8578] = 3'b110;
        rom_memory[8579] = 3'b110;
        rom_memory[8580] = 3'b110;
        rom_memory[8581] = 3'b110;
        rom_memory[8582] = 3'b110;
        rom_memory[8583] = 3'b110;
        rom_memory[8584] = 3'b110;
        rom_memory[8585] = 3'b110;
        rom_memory[8586] = 3'b110;
        rom_memory[8587] = 3'b110;
        rom_memory[8588] = 3'b110;
        rom_memory[8589] = 3'b110;
        rom_memory[8590] = 3'b110;
        rom_memory[8591] = 3'b110;
        rom_memory[8592] = 3'b110;
        rom_memory[8593] = 3'b110;
        rom_memory[8594] = 3'b110;
        rom_memory[8595] = 3'b110;
        rom_memory[8596] = 3'b110;
        rom_memory[8597] = 3'b110;
        rom_memory[8598] = 3'b110;
        rom_memory[8599] = 3'b110;
        rom_memory[8600] = 3'b110;
        rom_memory[8601] = 3'b110;
        rom_memory[8602] = 3'b110;
        rom_memory[8603] = 3'b110;
        rom_memory[8604] = 3'b110;
        rom_memory[8605] = 3'b110;
        rom_memory[8606] = 3'b110;
        rom_memory[8607] = 3'b110;
        rom_memory[8608] = 3'b110;
        rom_memory[8609] = 3'b110;
        rom_memory[8610] = 3'b110;
        rom_memory[8611] = 3'b110;
        rom_memory[8612] = 3'b110;
        rom_memory[8613] = 3'b110;
        rom_memory[8614] = 3'b110;
        rom_memory[8615] = 3'b110;
        rom_memory[8616] = 3'b110;
        rom_memory[8617] = 3'b110;
        rom_memory[8618] = 3'b110;
        rom_memory[8619] = 3'b110;
        rom_memory[8620] = 3'b110;
        rom_memory[8621] = 3'b110;
        rom_memory[8622] = 3'b110;
        rom_memory[8623] = 3'b110;
        rom_memory[8624] = 3'b110;
        rom_memory[8625] = 3'b110;
        rom_memory[8626] = 3'b110;
        rom_memory[8627] = 3'b110;
        rom_memory[8628] = 3'b110;
        rom_memory[8629] = 3'b110;
        rom_memory[8630] = 3'b110;
        rom_memory[8631] = 3'b110;
        rom_memory[8632] = 3'b110;
        rom_memory[8633] = 3'b110;
        rom_memory[8634] = 3'b110;
        rom_memory[8635] = 3'b110;
        rom_memory[8636] = 3'b110;
        rom_memory[8637] = 3'b110;
        rom_memory[8638] = 3'b110;
        rom_memory[8639] = 3'b110;
        rom_memory[8640] = 3'b110;
        rom_memory[8641] = 3'b110;
        rom_memory[8642] = 3'b110;
        rom_memory[8643] = 3'b110;
        rom_memory[8644] = 3'b110;
        rom_memory[8645] = 3'b110;
        rom_memory[8646] = 3'b110;
        rom_memory[8647] = 3'b110;
        rom_memory[8648] = 3'b110;
        rom_memory[8649] = 3'b110;
        rom_memory[8650] = 3'b110;
        rom_memory[8651] = 3'b110;
        rom_memory[8652] = 3'b110;
        rom_memory[8653] = 3'b110;
        rom_memory[8654] = 3'b110;
        rom_memory[8655] = 3'b110;
        rom_memory[8656] = 3'b110;
        rom_memory[8657] = 3'b110;
        rom_memory[8658] = 3'b110;
        rom_memory[8659] = 3'b110;
        rom_memory[8660] = 3'b110;
        rom_memory[8661] = 3'b110;
        rom_memory[8662] = 3'b110;
        rom_memory[8663] = 3'b110;
        rom_memory[8664] = 3'b110;
        rom_memory[8665] = 3'b110;
        rom_memory[8666] = 3'b110;
        rom_memory[8667] = 3'b110;
        rom_memory[8668] = 3'b110;
        rom_memory[8669] = 3'b110;
        rom_memory[8670] = 3'b110;
        rom_memory[8671] = 3'b110;
        rom_memory[8672] = 3'b110;
        rom_memory[8673] = 3'b110;
        rom_memory[8674] = 3'b110;
        rom_memory[8675] = 3'b110;
        rom_memory[8676] = 3'b110;
        rom_memory[8677] = 3'b110;
        rom_memory[8678] = 3'b110;
        rom_memory[8679] = 3'b110;
        rom_memory[8680] = 3'b110;
        rom_memory[8681] = 3'b110;
        rom_memory[8682] = 3'b110;
        rom_memory[8683] = 3'b110;
        rom_memory[8684] = 3'b110;
        rom_memory[8685] = 3'b111;
        rom_memory[8686] = 3'b000;
        rom_memory[8687] = 3'b000;
        rom_memory[8688] = 3'b000;
        rom_memory[8689] = 3'b000;
        rom_memory[8690] = 3'b000;
        rom_memory[8691] = 3'b000;
        rom_memory[8692] = 3'b000;
        rom_memory[8693] = 3'b000;
        rom_memory[8694] = 3'b000;
        rom_memory[8695] = 3'b000;
        rom_memory[8696] = 3'b000;
        rom_memory[8697] = 3'b000;
        rom_memory[8698] = 3'b000;
        rom_memory[8699] = 3'b000;
        rom_memory[8700] = 3'b000;
        rom_memory[8701] = 3'b000;
        rom_memory[8702] = 3'b000;
        rom_memory[8703] = 3'b000;
        rom_memory[8704] = 3'b001;
        rom_memory[8705] = 3'b000;
        rom_memory[8706] = 3'b000;
        rom_memory[8707] = 3'b000;
        rom_memory[8708] = 3'b000;
        rom_memory[8709] = 3'b000;
        rom_memory[8710] = 3'b000;
        rom_memory[8711] = 3'b000;
        rom_memory[8712] = 3'b000;
        rom_memory[8713] = 3'b000;
        rom_memory[8714] = 3'b000;
        rom_memory[8715] = 3'b000;
        rom_memory[8716] = 3'b000;
        rom_memory[8717] = 3'b000;
        rom_memory[8718] = 3'b000;
        rom_memory[8719] = 3'b000;
        rom_memory[8720] = 3'b000;
        rom_memory[8721] = 3'b000;
        rom_memory[8722] = 3'b000;
        rom_memory[8723] = 3'b010;
        rom_memory[8724] = 3'b000;
        rom_memory[8725] = 3'b010;
        rom_memory[8726] = 3'b011;
        rom_memory[8727] = 3'b011;
        rom_memory[8728] = 3'b011;
        rom_memory[8729] = 3'b011;
        rom_memory[8730] = 3'b011;
        rom_memory[8731] = 3'b011;
        rom_memory[8732] = 3'b011;
        rom_memory[8733] = 3'b001;
        rom_memory[8734] = 3'b111;
        rom_memory[8735] = 3'b110;
        rom_memory[8736] = 3'b110;
        rom_memory[8737] = 3'b110;
        rom_memory[8738] = 3'b110;
        rom_memory[8739] = 3'b110;
        rom_memory[8740] = 3'b110;
        rom_memory[8741] = 3'b110;
        rom_memory[8742] = 3'b110;
        rom_memory[8743] = 3'b110;
        rom_memory[8744] = 3'b110;
        rom_memory[8745] = 3'b110;
        rom_memory[8746] = 3'b110;
        rom_memory[8747] = 3'b110;
        rom_memory[8748] = 3'b110;
        rom_memory[8749] = 3'b110;
        rom_memory[8750] = 3'b110;
        rom_memory[8751] = 3'b110;
        rom_memory[8752] = 3'b110;
        rom_memory[8753] = 3'b110;
        rom_memory[8754] = 3'b110;
        rom_memory[8755] = 3'b110;
        rom_memory[8756] = 3'b110;
        rom_memory[8757] = 3'b110;
        rom_memory[8758] = 3'b110;
        rom_memory[8759] = 3'b110;
        rom_memory[8760] = 3'b110;
        rom_memory[8761] = 3'b110;
        rom_memory[8762] = 3'b110;
        rom_memory[8763] = 3'b110;
        rom_memory[8764] = 3'b110;
        rom_memory[8765] = 3'b110;
        rom_memory[8766] = 3'b110;
        rom_memory[8767] = 3'b110;
        rom_memory[8768] = 3'b110;
        rom_memory[8769] = 3'b110;
        rom_memory[8770] = 3'b110;
        rom_memory[8771] = 3'b110;
        rom_memory[8772] = 3'b110;
        rom_memory[8773] = 3'b110;
        rom_memory[8774] = 3'b110;
        rom_memory[8775] = 3'b110;
        rom_memory[8776] = 3'b110;
        rom_memory[8777] = 3'b110;
        rom_memory[8778] = 3'b110;
        rom_memory[8779] = 3'b110;
        rom_memory[8780] = 3'b110;
        rom_memory[8781] = 3'b110;
        rom_memory[8782] = 3'b110;
        rom_memory[8783] = 3'b110;
        rom_memory[8784] = 3'b110;
        rom_memory[8785] = 3'b110;
        rom_memory[8786] = 3'b110;
        rom_memory[8787] = 3'b110;
        rom_memory[8788] = 3'b110;
        rom_memory[8789] = 3'b110;
        rom_memory[8790] = 3'b110;
        rom_memory[8791] = 3'b110;
        rom_memory[8792] = 3'b110;
        rom_memory[8793] = 3'b110;
        rom_memory[8794] = 3'b110;
        rom_memory[8795] = 3'b110;
        rom_memory[8796] = 3'b110;
        rom_memory[8797] = 3'b110;
        rom_memory[8798] = 3'b110;
        rom_memory[8799] = 3'b110;
        rom_memory[8800] = 3'b110;
        rom_memory[8801] = 3'b110;
        rom_memory[8802] = 3'b110;
        rom_memory[8803] = 3'b110;
        rom_memory[8804] = 3'b110;
        rom_memory[8805] = 3'b110;
        rom_memory[8806] = 3'b110;
        rom_memory[8807] = 3'b110;
        rom_memory[8808] = 3'b110;
        rom_memory[8809] = 3'b110;
        rom_memory[8810] = 3'b110;
        rom_memory[8811] = 3'b110;
        rom_memory[8812] = 3'b110;
        rom_memory[8813] = 3'b110;
        rom_memory[8814] = 3'b110;
        rom_memory[8815] = 3'b110;
        rom_memory[8816] = 3'b110;
        rom_memory[8817] = 3'b110;
        rom_memory[8818] = 3'b110;
        rom_memory[8819] = 3'b110;
        rom_memory[8820] = 3'b110;
        rom_memory[8821] = 3'b110;
        rom_memory[8822] = 3'b110;
        rom_memory[8823] = 3'b110;
        rom_memory[8824] = 3'b110;
        rom_memory[8825] = 3'b110;
        rom_memory[8826] = 3'b110;
        rom_memory[8827] = 3'b110;
        rom_memory[8828] = 3'b110;
        rom_memory[8829] = 3'b110;
        rom_memory[8830] = 3'b110;
        rom_memory[8831] = 3'b110;
        rom_memory[8832] = 3'b110;
        rom_memory[8833] = 3'b110;
        rom_memory[8834] = 3'b110;
        rom_memory[8835] = 3'b110;
        rom_memory[8836] = 3'b110;
        rom_memory[8837] = 3'b110;
        rom_memory[8838] = 3'b110;
        rom_memory[8839] = 3'b110;
        rom_memory[8840] = 3'b110;
        rom_memory[8841] = 3'b110;
        rom_memory[8842] = 3'b110;
        rom_memory[8843] = 3'b110;
        rom_memory[8844] = 3'b110;
        rom_memory[8845] = 3'b110;
        rom_memory[8846] = 3'b110;
        rom_memory[8847] = 3'b110;
        rom_memory[8848] = 3'b110;
        rom_memory[8849] = 3'b110;
        rom_memory[8850] = 3'b110;
        rom_memory[8851] = 3'b110;
        rom_memory[8852] = 3'b110;
        rom_memory[8853] = 3'b110;
        rom_memory[8854] = 3'b110;
        rom_memory[8855] = 3'b110;
        rom_memory[8856] = 3'b110;
        rom_memory[8857] = 3'b110;
        rom_memory[8858] = 3'b110;
        rom_memory[8859] = 3'b110;
        rom_memory[8860] = 3'b110;
        rom_memory[8861] = 3'b110;
        rom_memory[8862] = 3'b110;
        rom_memory[8863] = 3'b110;
        rom_memory[8864] = 3'b110;
        rom_memory[8865] = 3'b110;
        rom_memory[8866] = 3'b110;
        rom_memory[8867] = 3'b110;
        rom_memory[8868] = 3'b110;
        rom_memory[8869] = 3'b110;
        rom_memory[8870] = 3'b110;
        rom_memory[8871] = 3'b110;
        rom_memory[8872] = 3'b110;
        rom_memory[8873] = 3'b110;
        rom_memory[8874] = 3'b110;
        rom_memory[8875] = 3'b110;
        rom_memory[8876] = 3'b110;
        rom_memory[8877] = 3'b110;
        rom_memory[8878] = 3'b110;
        rom_memory[8879] = 3'b110;
        rom_memory[8880] = 3'b110;
        rom_memory[8881] = 3'b110;
        rom_memory[8882] = 3'b110;
        rom_memory[8883] = 3'b110;
        rom_memory[8884] = 3'b110;
        rom_memory[8885] = 3'b110;
        rom_memory[8886] = 3'b110;
        rom_memory[8887] = 3'b110;
        rom_memory[8888] = 3'b110;
        rom_memory[8889] = 3'b110;
        rom_memory[8890] = 3'b110;
        rom_memory[8891] = 3'b110;
        rom_memory[8892] = 3'b110;
        rom_memory[8893] = 3'b110;
        rom_memory[8894] = 3'b110;
        rom_memory[8895] = 3'b110;
        rom_memory[8896] = 3'b110;
        rom_memory[8897] = 3'b110;
        rom_memory[8898] = 3'b110;
        rom_memory[8899] = 3'b110;
        rom_memory[8900] = 3'b110;
        rom_memory[8901] = 3'b110;
        rom_memory[8902] = 3'b110;
        rom_memory[8903] = 3'b110;
        rom_memory[8904] = 3'b110;
        rom_memory[8905] = 3'b110;
        rom_memory[8906] = 3'b110;
        rom_memory[8907] = 3'b110;
        rom_memory[8908] = 3'b110;
        rom_memory[8909] = 3'b110;
        rom_memory[8910] = 3'b110;
        rom_memory[8911] = 3'b110;
        rom_memory[8912] = 3'b110;
        rom_memory[8913] = 3'b110;
        rom_memory[8914] = 3'b110;
        rom_memory[8915] = 3'b110;
        rom_memory[8916] = 3'b110;
        rom_memory[8917] = 3'b110;
        rom_memory[8918] = 3'b110;
        rom_memory[8919] = 3'b110;
        rom_memory[8920] = 3'b110;
        rom_memory[8921] = 3'b110;
        rom_memory[8922] = 3'b110;
        rom_memory[8923] = 3'b110;
        rom_memory[8924] = 3'b110;
        rom_memory[8925] = 3'b111;
        rom_memory[8926] = 3'b110;
        rom_memory[8927] = 3'b000;
        rom_memory[8928] = 3'b000;
        rom_memory[8929] = 3'b000;
        rom_memory[8930] = 3'b000;
        rom_memory[8931] = 3'b000;
        rom_memory[8932] = 3'b000;
        rom_memory[8933] = 3'b000;
        rom_memory[8934] = 3'b000;
        rom_memory[8935] = 3'b000;
        rom_memory[8936] = 3'b000;
        rom_memory[8937] = 3'b000;
        rom_memory[8938] = 3'b000;
        rom_memory[8939] = 3'b000;
        rom_memory[8940] = 3'b000;
        rom_memory[8941] = 3'b000;
        rom_memory[8942] = 3'b000;
        rom_memory[8943] = 3'b000;
        rom_memory[8944] = 3'b000;
        rom_memory[8945] = 3'b000;
        rom_memory[8946] = 3'b000;
        rom_memory[8947] = 3'b000;
        rom_memory[8948] = 3'b000;
        rom_memory[8949] = 3'b000;
        rom_memory[8950] = 3'b000;
        rom_memory[8951] = 3'b000;
        rom_memory[8952] = 3'b000;
        rom_memory[8953] = 3'b000;
        rom_memory[8954] = 3'b000;
        rom_memory[8955] = 3'b000;
        rom_memory[8956] = 3'b000;
        rom_memory[8957] = 3'b000;
        rom_memory[8958] = 3'b000;
        rom_memory[8959] = 3'b000;
        rom_memory[8960] = 3'b000;
        rom_memory[8961] = 3'b000;
        rom_memory[8962] = 3'b011;
        rom_memory[8963] = 3'b010;
        rom_memory[8964] = 3'b010;
        rom_memory[8965] = 3'b011;
        rom_memory[8966] = 3'b000;
        rom_memory[8967] = 3'b011;
        rom_memory[8968] = 3'b011;
        rom_memory[8969] = 3'b011;
        rom_memory[8970] = 3'b011;
        rom_memory[8971] = 3'b001;
        rom_memory[8972] = 3'b011;
        rom_memory[8973] = 3'b011;
        rom_memory[8974] = 3'b000;
        rom_memory[8975] = 3'b111;
        rom_memory[8976] = 3'b110;
        rom_memory[8977] = 3'b110;
        rom_memory[8978] = 3'b110;
        rom_memory[8979] = 3'b110;
        rom_memory[8980] = 3'b110;
        rom_memory[8981] = 3'b110;
        rom_memory[8982] = 3'b110;
        rom_memory[8983] = 3'b110;
        rom_memory[8984] = 3'b110;
        rom_memory[8985] = 3'b110;
        rom_memory[8986] = 3'b110;
        rom_memory[8987] = 3'b110;
        rom_memory[8988] = 3'b110;
        rom_memory[8989] = 3'b110;
        rom_memory[8990] = 3'b110;
        rom_memory[8991] = 3'b110;
        rom_memory[8992] = 3'b110;
        rom_memory[8993] = 3'b110;
        rom_memory[8994] = 3'b110;
        rom_memory[8995] = 3'b110;
        rom_memory[8996] = 3'b110;
        rom_memory[8997] = 3'b110;
        rom_memory[8998] = 3'b110;
        rom_memory[8999] = 3'b110;
        rom_memory[9000] = 3'b110;
        rom_memory[9001] = 3'b110;
        rom_memory[9002] = 3'b110;
        rom_memory[9003] = 3'b110;
        rom_memory[9004] = 3'b110;
        rom_memory[9005] = 3'b110;
        rom_memory[9006] = 3'b110;
        rom_memory[9007] = 3'b110;
        rom_memory[9008] = 3'b110;
        rom_memory[9009] = 3'b110;
        rom_memory[9010] = 3'b110;
        rom_memory[9011] = 3'b110;
        rom_memory[9012] = 3'b110;
        rom_memory[9013] = 3'b110;
        rom_memory[9014] = 3'b110;
        rom_memory[9015] = 3'b110;
        rom_memory[9016] = 3'b110;
        rom_memory[9017] = 3'b110;
        rom_memory[9018] = 3'b110;
        rom_memory[9019] = 3'b110;
        rom_memory[9020] = 3'b110;
        rom_memory[9021] = 3'b110;
        rom_memory[9022] = 3'b110;
        rom_memory[9023] = 3'b110;
        rom_memory[9024] = 3'b110;
        rom_memory[9025] = 3'b110;
        rom_memory[9026] = 3'b110;
        rom_memory[9027] = 3'b110;
        rom_memory[9028] = 3'b110;
        rom_memory[9029] = 3'b110;
        rom_memory[9030] = 3'b110;
        rom_memory[9031] = 3'b110;
        rom_memory[9032] = 3'b110;
        rom_memory[9033] = 3'b110;
        rom_memory[9034] = 3'b110;
        rom_memory[9035] = 3'b110;
        rom_memory[9036] = 3'b110;
        rom_memory[9037] = 3'b110;
        rom_memory[9038] = 3'b110;
        rom_memory[9039] = 3'b110;
        rom_memory[9040] = 3'b110;
        rom_memory[9041] = 3'b110;
        rom_memory[9042] = 3'b110;
        rom_memory[9043] = 3'b110;
        rom_memory[9044] = 3'b110;
        rom_memory[9045] = 3'b110;
        rom_memory[9046] = 3'b110;
        rom_memory[9047] = 3'b110;
        rom_memory[9048] = 3'b110;
        rom_memory[9049] = 3'b110;
        rom_memory[9050] = 3'b110;
        rom_memory[9051] = 3'b110;
        rom_memory[9052] = 3'b110;
        rom_memory[9053] = 3'b110;
        rom_memory[9054] = 3'b110;
        rom_memory[9055] = 3'b110;
        rom_memory[9056] = 3'b110;
        rom_memory[9057] = 3'b110;
        rom_memory[9058] = 3'b110;
        rom_memory[9059] = 3'b110;
        rom_memory[9060] = 3'b110;
        rom_memory[9061] = 3'b110;
        rom_memory[9062] = 3'b110;
        rom_memory[9063] = 3'b110;
        rom_memory[9064] = 3'b110;
        rom_memory[9065] = 3'b110;
        rom_memory[9066] = 3'b110;
        rom_memory[9067] = 3'b110;
        rom_memory[9068] = 3'b110;
        rom_memory[9069] = 3'b110;
        rom_memory[9070] = 3'b110;
        rom_memory[9071] = 3'b110;
        rom_memory[9072] = 3'b110;
        rom_memory[9073] = 3'b110;
        rom_memory[9074] = 3'b110;
        rom_memory[9075] = 3'b110;
        rom_memory[9076] = 3'b110;
        rom_memory[9077] = 3'b110;
        rom_memory[9078] = 3'b110;
        rom_memory[9079] = 3'b110;
        rom_memory[9080] = 3'b110;
        rom_memory[9081] = 3'b110;
        rom_memory[9082] = 3'b110;
        rom_memory[9083] = 3'b110;
        rom_memory[9084] = 3'b110;
        rom_memory[9085] = 3'b110;
        rom_memory[9086] = 3'b110;
        rom_memory[9087] = 3'b110;
        rom_memory[9088] = 3'b110;
        rom_memory[9089] = 3'b110;
        rom_memory[9090] = 3'b110;
        rom_memory[9091] = 3'b110;
        rom_memory[9092] = 3'b110;
        rom_memory[9093] = 3'b110;
        rom_memory[9094] = 3'b110;
        rom_memory[9095] = 3'b110;
        rom_memory[9096] = 3'b110;
        rom_memory[9097] = 3'b110;
        rom_memory[9098] = 3'b110;
        rom_memory[9099] = 3'b110;
        rom_memory[9100] = 3'b110;
        rom_memory[9101] = 3'b110;
        rom_memory[9102] = 3'b110;
        rom_memory[9103] = 3'b110;
        rom_memory[9104] = 3'b110;
        rom_memory[9105] = 3'b110;
        rom_memory[9106] = 3'b110;
        rom_memory[9107] = 3'b110;
        rom_memory[9108] = 3'b110;
        rom_memory[9109] = 3'b110;
        rom_memory[9110] = 3'b110;
        rom_memory[9111] = 3'b110;
        rom_memory[9112] = 3'b110;
        rom_memory[9113] = 3'b110;
        rom_memory[9114] = 3'b110;
        rom_memory[9115] = 3'b110;
        rom_memory[9116] = 3'b110;
        rom_memory[9117] = 3'b110;
        rom_memory[9118] = 3'b110;
        rom_memory[9119] = 3'b110;
        rom_memory[9120] = 3'b110;
        rom_memory[9121] = 3'b110;
        rom_memory[9122] = 3'b110;
        rom_memory[9123] = 3'b110;
        rom_memory[9124] = 3'b110;
        rom_memory[9125] = 3'b110;
        rom_memory[9126] = 3'b110;
        rom_memory[9127] = 3'b110;
        rom_memory[9128] = 3'b110;
        rom_memory[9129] = 3'b110;
        rom_memory[9130] = 3'b110;
        rom_memory[9131] = 3'b110;
        rom_memory[9132] = 3'b110;
        rom_memory[9133] = 3'b110;
        rom_memory[9134] = 3'b110;
        rom_memory[9135] = 3'b110;
        rom_memory[9136] = 3'b110;
        rom_memory[9137] = 3'b110;
        rom_memory[9138] = 3'b110;
        rom_memory[9139] = 3'b110;
        rom_memory[9140] = 3'b110;
        rom_memory[9141] = 3'b110;
        rom_memory[9142] = 3'b110;
        rom_memory[9143] = 3'b110;
        rom_memory[9144] = 3'b110;
        rom_memory[9145] = 3'b110;
        rom_memory[9146] = 3'b110;
        rom_memory[9147] = 3'b110;
        rom_memory[9148] = 3'b110;
        rom_memory[9149] = 3'b110;
        rom_memory[9150] = 3'b110;
        rom_memory[9151] = 3'b110;
        rom_memory[9152] = 3'b110;
        rom_memory[9153] = 3'b110;
        rom_memory[9154] = 3'b110;
        rom_memory[9155] = 3'b110;
        rom_memory[9156] = 3'b110;
        rom_memory[9157] = 3'b110;
        rom_memory[9158] = 3'b110;
        rom_memory[9159] = 3'b110;
        rom_memory[9160] = 3'b110;
        rom_memory[9161] = 3'b110;
        rom_memory[9162] = 3'b110;
        rom_memory[9163] = 3'b110;
        rom_memory[9164] = 3'b110;
        rom_memory[9165] = 3'b111;
        rom_memory[9166] = 3'b110;
        rom_memory[9167] = 3'b000;
        rom_memory[9168] = 3'b000;
        rom_memory[9169] = 3'b000;
        rom_memory[9170] = 3'b000;
        rom_memory[9171] = 3'b000;
        rom_memory[9172] = 3'b000;
        rom_memory[9173] = 3'b000;
        rom_memory[9174] = 3'b000;
        rom_memory[9175] = 3'b000;
        rom_memory[9176] = 3'b000;
        rom_memory[9177] = 3'b000;
        rom_memory[9178] = 3'b000;
        rom_memory[9179] = 3'b000;
        rom_memory[9180] = 3'b000;
        rom_memory[9181] = 3'b000;
        rom_memory[9182] = 3'b000;
        rom_memory[9183] = 3'b000;
        rom_memory[9184] = 3'b000;
        rom_memory[9185] = 3'b000;
        rom_memory[9186] = 3'b000;
        rom_memory[9187] = 3'b000;
        rom_memory[9188] = 3'b000;
        rom_memory[9189] = 3'b000;
        rom_memory[9190] = 3'b000;
        rom_memory[9191] = 3'b000;
        rom_memory[9192] = 3'b000;
        rom_memory[9193] = 3'b000;
        rom_memory[9194] = 3'b000;
        rom_memory[9195] = 3'b000;
        rom_memory[9196] = 3'b000;
        rom_memory[9197] = 3'b000;
        rom_memory[9198] = 3'b000;
        rom_memory[9199] = 3'b000;
        rom_memory[9200] = 3'b000;
        rom_memory[9201] = 3'b000;
        rom_memory[9202] = 3'b010;
        rom_memory[9203] = 3'b010;
        rom_memory[9204] = 3'b010;
        rom_memory[9205] = 3'b011;
        rom_memory[9206] = 3'b011;
        rom_memory[9207] = 3'b011;
        rom_memory[9208] = 3'b011;
        rom_memory[9209] = 3'b011;
        rom_memory[9210] = 3'b011;
        rom_memory[9211] = 3'b011;
        rom_memory[9212] = 3'b011;
        rom_memory[9213] = 3'b011;
        rom_memory[9214] = 3'b111;
        rom_memory[9215] = 3'b111;
        rom_memory[9216] = 3'b111;
        rom_memory[9217] = 3'b110;
        rom_memory[9218] = 3'b111;
        rom_memory[9219] = 3'b110;
        rom_memory[9220] = 3'b110;
        rom_memory[9221] = 3'b110;
        rom_memory[9222] = 3'b110;
        rom_memory[9223] = 3'b110;
        rom_memory[9224] = 3'b111;
        rom_memory[9225] = 3'b110;
        rom_memory[9226] = 3'b110;
        rom_memory[9227] = 3'b110;
        rom_memory[9228] = 3'b110;
        rom_memory[9229] = 3'b110;
        rom_memory[9230] = 3'b110;
        rom_memory[9231] = 3'b110;
        rom_memory[9232] = 3'b110;
        rom_memory[9233] = 3'b110;
        rom_memory[9234] = 3'b110;
        rom_memory[9235] = 3'b110;
        rom_memory[9236] = 3'b110;
        rom_memory[9237] = 3'b110;
        rom_memory[9238] = 3'b110;
        rom_memory[9239] = 3'b110;
        rom_memory[9240] = 3'b110;
        rom_memory[9241] = 3'b110;
        rom_memory[9242] = 3'b110;
        rom_memory[9243] = 3'b110;
        rom_memory[9244] = 3'b110;
        rom_memory[9245] = 3'b110;
        rom_memory[9246] = 3'b110;
        rom_memory[9247] = 3'b110;
        rom_memory[9248] = 3'b110;
        rom_memory[9249] = 3'b110;
        rom_memory[9250] = 3'b110;
        rom_memory[9251] = 3'b110;
        rom_memory[9252] = 3'b110;
        rom_memory[9253] = 3'b110;
        rom_memory[9254] = 3'b110;
        rom_memory[9255] = 3'b110;
        rom_memory[9256] = 3'b110;
        rom_memory[9257] = 3'b110;
        rom_memory[9258] = 3'b110;
        rom_memory[9259] = 3'b110;
        rom_memory[9260] = 3'b110;
        rom_memory[9261] = 3'b110;
        rom_memory[9262] = 3'b110;
        rom_memory[9263] = 3'b110;
        rom_memory[9264] = 3'b110;
        rom_memory[9265] = 3'b110;
        rom_memory[9266] = 3'b110;
        rom_memory[9267] = 3'b110;
        rom_memory[9268] = 3'b110;
        rom_memory[9269] = 3'b110;
        rom_memory[9270] = 3'b110;
        rom_memory[9271] = 3'b110;
        rom_memory[9272] = 3'b110;
        rom_memory[9273] = 3'b110;
        rom_memory[9274] = 3'b110;
        rom_memory[9275] = 3'b110;
        rom_memory[9276] = 3'b110;
        rom_memory[9277] = 3'b110;
        rom_memory[9278] = 3'b110;
        rom_memory[9279] = 3'b110;
        rom_memory[9280] = 3'b110;
        rom_memory[9281] = 3'b110;
        rom_memory[9282] = 3'b110;
        rom_memory[9283] = 3'b110;
        rom_memory[9284] = 3'b110;
        rom_memory[9285] = 3'b110;
        rom_memory[9286] = 3'b110;
        rom_memory[9287] = 3'b110;
        rom_memory[9288] = 3'b110;
        rom_memory[9289] = 3'b110;
        rom_memory[9290] = 3'b110;
        rom_memory[9291] = 3'b110;
        rom_memory[9292] = 3'b110;
        rom_memory[9293] = 3'b110;
        rom_memory[9294] = 3'b110;
        rom_memory[9295] = 3'b110;
        rom_memory[9296] = 3'b110;
        rom_memory[9297] = 3'b110;
        rom_memory[9298] = 3'b110;
        rom_memory[9299] = 3'b110;
        rom_memory[9300] = 3'b110;
        rom_memory[9301] = 3'b110;
        rom_memory[9302] = 3'b110;
        rom_memory[9303] = 3'b110;
        rom_memory[9304] = 3'b110;
        rom_memory[9305] = 3'b110;
        rom_memory[9306] = 3'b110;
        rom_memory[9307] = 3'b110;
        rom_memory[9308] = 3'b110;
        rom_memory[9309] = 3'b110;
        rom_memory[9310] = 3'b110;
        rom_memory[9311] = 3'b110;
        rom_memory[9312] = 3'b110;
        rom_memory[9313] = 3'b110;
        rom_memory[9314] = 3'b110;
        rom_memory[9315] = 3'b110;
        rom_memory[9316] = 3'b110;
        rom_memory[9317] = 3'b110;
        rom_memory[9318] = 3'b110;
        rom_memory[9319] = 3'b110;
        rom_memory[9320] = 3'b110;
        rom_memory[9321] = 3'b110;
        rom_memory[9322] = 3'b110;
        rom_memory[9323] = 3'b110;
        rom_memory[9324] = 3'b110;
        rom_memory[9325] = 3'b110;
        rom_memory[9326] = 3'b110;
        rom_memory[9327] = 3'b110;
        rom_memory[9328] = 3'b110;
        rom_memory[9329] = 3'b110;
        rom_memory[9330] = 3'b110;
        rom_memory[9331] = 3'b110;
        rom_memory[9332] = 3'b110;
        rom_memory[9333] = 3'b110;
        rom_memory[9334] = 3'b110;
        rom_memory[9335] = 3'b110;
        rom_memory[9336] = 3'b110;
        rom_memory[9337] = 3'b110;
        rom_memory[9338] = 3'b110;
        rom_memory[9339] = 3'b110;
        rom_memory[9340] = 3'b110;
        rom_memory[9341] = 3'b110;
        rom_memory[9342] = 3'b110;
        rom_memory[9343] = 3'b110;
        rom_memory[9344] = 3'b110;
        rom_memory[9345] = 3'b110;
        rom_memory[9346] = 3'b110;
        rom_memory[9347] = 3'b110;
        rom_memory[9348] = 3'b110;
        rom_memory[9349] = 3'b110;
        rom_memory[9350] = 3'b110;
        rom_memory[9351] = 3'b110;
        rom_memory[9352] = 3'b110;
        rom_memory[9353] = 3'b110;
        rom_memory[9354] = 3'b110;
        rom_memory[9355] = 3'b110;
        rom_memory[9356] = 3'b110;
        rom_memory[9357] = 3'b110;
        rom_memory[9358] = 3'b110;
        rom_memory[9359] = 3'b110;
        rom_memory[9360] = 3'b110;
        rom_memory[9361] = 3'b110;
        rom_memory[9362] = 3'b110;
        rom_memory[9363] = 3'b110;
        rom_memory[9364] = 3'b110;
        rom_memory[9365] = 3'b110;
        rom_memory[9366] = 3'b110;
        rom_memory[9367] = 3'b110;
        rom_memory[9368] = 3'b110;
        rom_memory[9369] = 3'b110;
        rom_memory[9370] = 3'b110;
        rom_memory[9371] = 3'b110;
        rom_memory[9372] = 3'b110;
        rom_memory[9373] = 3'b110;
        rom_memory[9374] = 3'b110;
        rom_memory[9375] = 3'b110;
        rom_memory[9376] = 3'b110;
        rom_memory[9377] = 3'b110;
        rom_memory[9378] = 3'b110;
        rom_memory[9379] = 3'b110;
        rom_memory[9380] = 3'b110;
        rom_memory[9381] = 3'b110;
        rom_memory[9382] = 3'b110;
        rom_memory[9383] = 3'b110;
        rom_memory[9384] = 3'b110;
        rom_memory[9385] = 3'b110;
        rom_memory[9386] = 3'b110;
        rom_memory[9387] = 3'b110;
        rom_memory[9388] = 3'b110;
        rom_memory[9389] = 3'b110;
        rom_memory[9390] = 3'b110;
        rom_memory[9391] = 3'b110;
        rom_memory[9392] = 3'b110;
        rom_memory[9393] = 3'b110;
        rom_memory[9394] = 3'b110;
        rom_memory[9395] = 3'b110;
        rom_memory[9396] = 3'b110;
        rom_memory[9397] = 3'b110;
        rom_memory[9398] = 3'b110;
        rom_memory[9399] = 3'b110;
        rom_memory[9400] = 3'b110;
        rom_memory[9401] = 3'b110;
        rom_memory[9402] = 3'b110;
        rom_memory[9403] = 3'b110;
        rom_memory[9404] = 3'b110;
        rom_memory[9405] = 3'b110;
        rom_memory[9406] = 3'b111;
        rom_memory[9407] = 3'b000;
        rom_memory[9408] = 3'b000;
        rom_memory[9409] = 3'b000;
        rom_memory[9410] = 3'b000;
        rom_memory[9411] = 3'b000;
        rom_memory[9412] = 3'b000;
        rom_memory[9413] = 3'b000;
        rom_memory[9414] = 3'b000;
        rom_memory[9415] = 3'b000;
        rom_memory[9416] = 3'b000;
        rom_memory[9417] = 3'b000;
        rom_memory[9418] = 3'b000;
        rom_memory[9419] = 3'b000;
        rom_memory[9420] = 3'b000;
        rom_memory[9421] = 3'b000;
        rom_memory[9422] = 3'b000;
        rom_memory[9423] = 3'b000;
        rom_memory[9424] = 3'b000;
        rom_memory[9425] = 3'b000;
        rom_memory[9426] = 3'b000;
        rom_memory[9427] = 3'b000;
        rom_memory[9428] = 3'b000;
        rom_memory[9429] = 3'b000;
        rom_memory[9430] = 3'b000;
        rom_memory[9431] = 3'b000;
        rom_memory[9432] = 3'b000;
        rom_memory[9433] = 3'b000;
        rom_memory[9434] = 3'b000;
        rom_memory[9435] = 3'b000;
        rom_memory[9436] = 3'b000;
        rom_memory[9437] = 3'b000;
        rom_memory[9438] = 3'b000;
        rom_memory[9439] = 3'b000;
        rom_memory[9440] = 3'b000;
        rom_memory[9441] = 3'b000;
        rom_memory[9442] = 3'b000;
        rom_memory[9443] = 3'b000;
        rom_memory[9444] = 3'b000;
        rom_memory[9445] = 3'b011;
        rom_memory[9446] = 3'b011;
        rom_memory[9447] = 3'b011;
        rom_memory[9448] = 3'b011;
        rom_memory[9449] = 3'b011;
        rom_memory[9450] = 3'b011;
        rom_memory[9451] = 3'b011;
        rom_memory[9452] = 3'b011;
        rom_memory[9453] = 3'b011;
        rom_memory[9454] = 3'b011;
        rom_memory[9455] = 3'b111;
        rom_memory[9456] = 3'b111;
        rom_memory[9457] = 3'b110;
        rom_memory[9458] = 3'b111;
        rom_memory[9459] = 3'b110;
        rom_memory[9460] = 3'b110;
        rom_memory[9461] = 3'b110;
        rom_memory[9462] = 3'b110;
        rom_memory[9463] = 3'b110;
        rom_memory[9464] = 3'b110;
        rom_memory[9465] = 3'b110;
        rom_memory[9466] = 3'b110;
        rom_memory[9467] = 3'b110;
        rom_memory[9468] = 3'b110;
        rom_memory[9469] = 3'b110;
        rom_memory[9470] = 3'b110;
        rom_memory[9471] = 3'b110;
        rom_memory[9472] = 3'b110;
        rom_memory[9473] = 3'b110;
        rom_memory[9474] = 3'b110;
        rom_memory[9475] = 3'b110;
        rom_memory[9476] = 3'b110;
        rom_memory[9477] = 3'b110;
        rom_memory[9478] = 3'b110;
        rom_memory[9479] = 3'b110;
        rom_memory[9480] = 3'b110;
        rom_memory[9481] = 3'b110;
        rom_memory[9482] = 3'b110;
        rom_memory[9483] = 3'b110;
        rom_memory[9484] = 3'b110;
        rom_memory[9485] = 3'b110;
        rom_memory[9486] = 3'b110;
        rom_memory[9487] = 3'b110;
        rom_memory[9488] = 3'b110;
        rom_memory[9489] = 3'b110;
        rom_memory[9490] = 3'b110;
        rom_memory[9491] = 3'b110;
        rom_memory[9492] = 3'b110;
        rom_memory[9493] = 3'b110;
        rom_memory[9494] = 3'b110;
        rom_memory[9495] = 3'b110;
        rom_memory[9496] = 3'b110;
        rom_memory[9497] = 3'b110;
        rom_memory[9498] = 3'b110;
        rom_memory[9499] = 3'b110;
        rom_memory[9500] = 3'b110;
        rom_memory[9501] = 3'b110;
        rom_memory[9502] = 3'b110;
        rom_memory[9503] = 3'b110;
        rom_memory[9504] = 3'b110;
        rom_memory[9505] = 3'b110;
        rom_memory[9506] = 3'b110;
        rom_memory[9507] = 3'b110;
        rom_memory[9508] = 3'b110;
        rom_memory[9509] = 3'b110;
        rom_memory[9510] = 3'b110;
        rom_memory[9511] = 3'b110;
        rom_memory[9512] = 3'b110;
        rom_memory[9513] = 3'b110;
        rom_memory[9514] = 3'b110;
        rom_memory[9515] = 3'b110;
        rom_memory[9516] = 3'b110;
        rom_memory[9517] = 3'b110;
        rom_memory[9518] = 3'b110;
        rom_memory[9519] = 3'b110;
        rom_memory[9520] = 3'b110;
        rom_memory[9521] = 3'b110;
        rom_memory[9522] = 3'b110;
        rom_memory[9523] = 3'b110;
        rom_memory[9524] = 3'b110;
        rom_memory[9525] = 3'b110;
        rom_memory[9526] = 3'b110;
        rom_memory[9527] = 3'b110;
        rom_memory[9528] = 3'b110;
        rom_memory[9529] = 3'b110;
        rom_memory[9530] = 3'b110;
        rom_memory[9531] = 3'b110;
        rom_memory[9532] = 3'b110;
        rom_memory[9533] = 3'b110;
        rom_memory[9534] = 3'b110;
        rom_memory[9535] = 3'b110;
        rom_memory[9536] = 3'b110;
        rom_memory[9537] = 3'b110;
        rom_memory[9538] = 3'b110;
        rom_memory[9539] = 3'b110;
        rom_memory[9540] = 3'b110;
        rom_memory[9541] = 3'b110;
        rom_memory[9542] = 3'b110;
        rom_memory[9543] = 3'b110;
        rom_memory[9544] = 3'b110;
        rom_memory[9545] = 3'b110;
        rom_memory[9546] = 3'b110;
        rom_memory[9547] = 3'b110;
        rom_memory[9548] = 3'b110;
        rom_memory[9549] = 3'b110;
        rom_memory[9550] = 3'b110;
        rom_memory[9551] = 3'b110;
        rom_memory[9552] = 3'b110;
        rom_memory[9553] = 3'b110;
        rom_memory[9554] = 3'b110;
        rom_memory[9555] = 3'b110;
        rom_memory[9556] = 3'b110;
        rom_memory[9557] = 3'b110;
        rom_memory[9558] = 3'b110;
        rom_memory[9559] = 3'b110;
        rom_memory[9560] = 3'b110;
        rom_memory[9561] = 3'b110;
        rom_memory[9562] = 3'b110;
        rom_memory[9563] = 3'b110;
        rom_memory[9564] = 3'b110;
        rom_memory[9565] = 3'b110;
        rom_memory[9566] = 3'b110;
        rom_memory[9567] = 3'b110;
        rom_memory[9568] = 3'b110;
        rom_memory[9569] = 3'b110;
        rom_memory[9570] = 3'b110;
        rom_memory[9571] = 3'b110;
        rom_memory[9572] = 3'b110;
        rom_memory[9573] = 3'b110;
        rom_memory[9574] = 3'b110;
        rom_memory[9575] = 3'b110;
        rom_memory[9576] = 3'b110;
        rom_memory[9577] = 3'b110;
        rom_memory[9578] = 3'b110;
        rom_memory[9579] = 3'b110;
        rom_memory[9580] = 3'b110;
        rom_memory[9581] = 3'b110;
        rom_memory[9582] = 3'b110;
        rom_memory[9583] = 3'b110;
        rom_memory[9584] = 3'b110;
        rom_memory[9585] = 3'b110;
        rom_memory[9586] = 3'b110;
        rom_memory[9587] = 3'b110;
        rom_memory[9588] = 3'b110;
        rom_memory[9589] = 3'b110;
        rom_memory[9590] = 3'b110;
        rom_memory[9591] = 3'b110;
        rom_memory[9592] = 3'b110;
        rom_memory[9593] = 3'b110;
        rom_memory[9594] = 3'b110;
        rom_memory[9595] = 3'b110;
        rom_memory[9596] = 3'b110;
        rom_memory[9597] = 3'b110;
        rom_memory[9598] = 3'b110;
        rom_memory[9599] = 3'b110;
        rom_memory[9600] = 3'b110;
        rom_memory[9601] = 3'b110;
        rom_memory[9602] = 3'b110;
        rom_memory[9603] = 3'b110;
        rom_memory[9604] = 3'b110;
        rom_memory[9605] = 3'b110;
        rom_memory[9606] = 3'b110;
        rom_memory[9607] = 3'b110;
        rom_memory[9608] = 3'b110;
        rom_memory[9609] = 3'b110;
        rom_memory[9610] = 3'b110;
        rom_memory[9611] = 3'b110;
        rom_memory[9612] = 3'b110;
        rom_memory[9613] = 3'b110;
        rom_memory[9614] = 3'b110;
        rom_memory[9615] = 3'b110;
        rom_memory[9616] = 3'b110;
        rom_memory[9617] = 3'b110;
        rom_memory[9618] = 3'b110;
        rom_memory[9619] = 3'b110;
        rom_memory[9620] = 3'b110;
        rom_memory[9621] = 3'b110;
        rom_memory[9622] = 3'b110;
        rom_memory[9623] = 3'b110;
        rom_memory[9624] = 3'b110;
        rom_memory[9625] = 3'b110;
        rom_memory[9626] = 3'b110;
        rom_memory[9627] = 3'b110;
        rom_memory[9628] = 3'b110;
        rom_memory[9629] = 3'b110;
        rom_memory[9630] = 3'b110;
        rom_memory[9631] = 3'b110;
        rom_memory[9632] = 3'b110;
        rom_memory[9633] = 3'b110;
        rom_memory[9634] = 3'b110;
        rom_memory[9635] = 3'b110;
        rom_memory[9636] = 3'b110;
        rom_memory[9637] = 3'b110;
        rom_memory[9638] = 3'b110;
        rom_memory[9639] = 3'b110;
        rom_memory[9640] = 3'b110;
        rom_memory[9641] = 3'b110;
        rom_memory[9642] = 3'b110;
        rom_memory[9643] = 3'b110;
        rom_memory[9644] = 3'b110;
        rom_memory[9645] = 3'b110;
        rom_memory[9646] = 3'b111;
        rom_memory[9647] = 3'b110;
        rom_memory[9648] = 3'b000;
        rom_memory[9649] = 3'b000;
        rom_memory[9650] = 3'b000;
        rom_memory[9651] = 3'b000;
        rom_memory[9652] = 3'b000;
        rom_memory[9653] = 3'b000;
        rom_memory[9654] = 3'b000;
        rom_memory[9655] = 3'b000;
        rom_memory[9656] = 3'b000;
        rom_memory[9657] = 3'b000;
        rom_memory[9658] = 3'b000;
        rom_memory[9659] = 3'b000;
        rom_memory[9660] = 3'b000;
        rom_memory[9661] = 3'b000;
        rom_memory[9662] = 3'b000;
        rom_memory[9663] = 3'b000;
        rom_memory[9664] = 3'b000;
        rom_memory[9665] = 3'b000;
        rom_memory[9666] = 3'b000;
        rom_memory[9667] = 3'b000;
        rom_memory[9668] = 3'b000;
        rom_memory[9669] = 3'b000;
        rom_memory[9670] = 3'b000;
        rom_memory[9671] = 3'b000;
        rom_memory[9672] = 3'b000;
        rom_memory[9673] = 3'b000;
        rom_memory[9674] = 3'b000;
        rom_memory[9675] = 3'b000;
        rom_memory[9676] = 3'b000;
        rom_memory[9677] = 3'b000;
        rom_memory[9678] = 3'b000;
        rom_memory[9679] = 3'b000;
        rom_memory[9680] = 3'b000;
        rom_memory[9681] = 3'b000;
        rom_memory[9682] = 3'b000;
        rom_memory[9683] = 3'b000;
        rom_memory[9684] = 3'b000;
        rom_memory[9685] = 3'b010;
        rom_memory[9686] = 3'b011;
        rom_memory[9687] = 3'b011;
        rom_memory[9688] = 3'b000;
        rom_memory[9689] = 3'b011;
        rom_memory[9690] = 3'b011;
        rom_memory[9691] = 3'b011;
        rom_memory[9692] = 3'b011;
        rom_memory[9693] = 3'b011;
        rom_memory[9694] = 3'b011;
        rom_memory[9695] = 3'b011;
        rom_memory[9696] = 3'b111;
        rom_memory[9697] = 3'b111;
        rom_memory[9698] = 3'b110;
        rom_memory[9699] = 3'b110;
        rom_memory[9700] = 3'b110;
        rom_memory[9701] = 3'b110;
        rom_memory[9702] = 3'b110;
        rom_memory[9703] = 3'b110;
        rom_memory[9704] = 3'b110;
        rom_memory[9705] = 3'b110;
        rom_memory[9706] = 3'b110;
        rom_memory[9707] = 3'b110;
        rom_memory[9708] = 3'b110;
        rom_memory[9709] = 3'b110;
        rom_memory[9710] = 3'b110;
        rom_memory[9711] = 3'b110;
        rom_memory[9712] = 3'b110;
        rom_memory[9713] = 3'b110;
        rom_memory[9714] = 3'b110;
        rom_memory[9715] = 3'b110;
        rom_memory[9716] = 3'b110;
        rom_memory[9717] = 3'b110;
        rom_memory[9718] = 3'b110;
        rom_memory[9719] = 3'b110;
        rom_memory[9720] = 3'b110;
        rom_memory[9721] = 3'b110;
        rom_memory[9722] = 3'b110;
        rom_memory[9723] = 3'b110;
        rom_memory[9724] = 3'b110;
        rom_memory[9725] = 3'b110;
        rom_memory[9726] = 3'b110;
        rom_memory[9727] = 3'b110;
        rom_memory[9728] = 3'b110;
        rom_memory[9729] = 3'b110;
        rom_memory[9730] = 3'b110;
        rom_memory[9731] = 3'b110;
        rom_memory[9732] = 3'b110;
        rom_memory[9733] = 3'b110;
        rom_memory[9734] = 3'b110;
        rom_memory[9735] = 3'b110;
        rom_memory[9736] = 3'b110;
        rom_memory[9737] = 3'b110;
        rom_memory[9738] = 3'b110;
        rom_memory[9739] = 3'b110;
        rom_memory[9740] = 3'b110;
        rom_memory[9741] = 3'b110;
        rom_memory[9742] = 3'b110;
        rom_memory[9743] = 3'b110;
        rom_memory[9744] = 3'b110;
        rom_memory[9745] = 3'b110;
        rom_memory[9746] = 3'b110;
        rom_memory[9747] = 3'b110;
        rom_memory[9748] = 3'b110;
        rom_memory[9749] = 3'b110;
        rom_memory[9750] = 3'b110;
        rom_memory[9751] = 3'b110;
        rom_memory[9752] = 3'b110;
        rom_memory[9753] = 3'b110;
        rom_memory[9754] = 3'b110;
        rom_memory[9755] = 3'b110;
        rom_memory[9756] = 3'b110;
        rom_memory[9757] = 3'b110;
        rom_memory[9758] = 3'b110;
        rom_memory[9759] = 3'b110;
        rom_memory[9760] = 3'b110;
        rom_memory[9761] = 3'b110;
        rom_memory[9762] = 3'b110;
        rom_memory[9763] = 3'b110;
        rom_memory[9764] = 3'b110;
        rom_memory[9765] = 3'b110;
        rom_memory[9766] = 3'b110;
        rom_memory[9767] = 3'b110;
        rom_memory[9768] = 3'b110;
        rom_memory[9769] = 3'b110;
        rom_memory[9770] = 3'b110;
        rom_memory[9771] = 3'b110;
        rom_memory[9772] = 3'b110;
        rom_memory[9773] = 3'b110;
        rom_memory[9774] = 3'b110;
        rom_memory[9775] = 3'b110;
        rom_memory[9776] = 3'b110;
        rom_memory[9777] = 3'b110;
        rom_memory[9778] = 3'b110;
        rom_memory[9779] = 3'b110;
        rom_memory[9780] = 3'b110;
        rom_memory[9781] = 3'b110;
        rom_memory[9782] = 3'b110;
        rom_memory[9783] = 3'b110;
        rom_memory[9784] = 3'b110;
        rom_memory[9785] = 3'b110;
        rom_memory[9786] = 3'b110;
        rom_memory[9787] = 3'b110;
        rom_memory[9788] = 3'b110;
        rom_memory[9789] = 3'b110;
        rom_memory[9790] = 3'b110;
        rom_memory[9791] = 3'b110;
        rom_memory[9792] = 3'b110;
        rom_memory[9793] = 3'b110;
        rom_memory[9794] = 3'b110;
        rom_memory[9795] = 3'b110;
        rom_memory[9796] = 3'b110;
        rom_memory[9797] = 3'b110;
        rom_memory[9798] = 3'b110;
        rom_memory[9799] = 3'b110;
        rom_memory[9800] = 3'b110;
        rom_memory[9801] = 3'b110;
        rom_memory[9802] = 3'b110;
        rom_memory[9803] = 3'b110;
        rom_memory[9804] = 3'b110;
        rom_memory[9805] = 3'b110;
        rom_memory[9806] = 3'b110;
        rom_memory[9807] = 3'b110;
        rom_memory[9808] = 3'b110;
        rom_memory[9809] = 3'b110;
        rom_memory[9810] = 3'b110;
        rom_memory[9811] = 3'b110;
        rom_memory[9812] = 3'b110;
        rom_memory[9813] = 3'b110;
        rom_memory[9814] = 3'b110;
        rom_memory[9815] = 3'b110;
        rom_memory[9816] = 3'b110;
        rom_memory[9817] = 3'b110;
        rom_memory[9818] = 3'b110;
        rom_memory[9819] = 3'b110;
        rom_memory[9820] = 3'b110;
        rom_memory[9821] = 3'b110;
        rom_memory[9822] = 3'b110;
        rom_memory[9823] = 3'b110;
        rom_memory[9824] = 3'b110;
        rom_memory[9825] = 3'b110;
        rom_memory[9826] = 3'b110;
        rom_memory[9827] = 3'b110;
        rom_memory[9828] = 3'b110;
        rom_memory[9829] = 3'b110;
        rom_memory[9830] = 3'b110;
        rom_memory[9831] = 3'b110;
        rom_memory[9832] = 3'b110;
        rom_memory[9833] = 3'b110;
        rom_memory[9834] = 3'b110;
        rom_memory[9835] = 3'b110;
        rom_memory[9836] = 3'b110;
        rom_memory[9837] = 3'b110;
        rom_memory[9838] = 3'b110;
        rom_memory[9839] = 3'b110;
        rom_memory[9840] = 3'b110;
        rom_memory[9841] = 3'b110;
        rom_memory[9842] = 3'b110;
        rom_memory[9843] = 3'b110;
        rom_memory[9844] = 3'b110;
        rom_memory[9845] = 3'b110;
        rom_memory[9846] = 3'b110;
        rom_memory[9847] = 3'b110;
        rom_memory[9848] = 3'b110;
        rom_memory[9849] = 3'b110;
        rom_memory[9850] = 3'b110;
        rom_memory[9851] = 3'b110;
        rom_memory[9852] = 3'b110;
        rom_memory[9853] = 3'b110;
        rom_memory[9854] = 3'b110;
        rom_memory[9855] = 3'b110;
        rom_memory[9856] = 3'b110;
        rom_memory[9857] = 3'b110;
        rom_memory[9858] = 3'b110;
        rom_memory[9859] = 3'b110;
        rom_memory[9860] = 3'b110;
        rom_memory[9861] = 3'b110;
        rom_memory[9862] = 3'b110;
        rom_memory[9863] = 3'b110;
        rom_memory[9864] = 3'b110;
        rom_memory[9865] = 3'b110;
        rom_memory[9866] = 3'b110;
        rom_memory[9867] = 3'b110;
        rom_memory[9868] = 3'b110;
        rom_memory[9869] = 3'b110;
        rom_memory[9870] = 3'b110;
        rom_memory[9871] = 3'b110;
        rom_memory[9872] = 3'b110;
        rom_memory[9873] = 3'b110;
        rom_memory[9874] = 3'b110;
        rom_memory[9875] = 3'b110;
        rom_memory[9876] = 3'b110;
        rom_memory[9877] = 3'b110;
        rom_memory[9878] = 3'b110;
        rom_memory[9879] = 3'b110;
        rom_memory[9880] = 3'b110;
        rom_memory[9881] = 3'b110;
        rom_memory[9882] = 3'b110;
        rom_memory[9883] = 3'b110;
        rom_memory[9884] = 3'b110;
        rom_memory[9885] = 3'b111;
        rom_memory[9886] = 3'b111;
        rom_memory[9887] = 3'b110;
        rom_memory[9888] = 3'b000;
        rom_memory[9889] = 3'b000;
        rom_memory[9890] = 3'b000;
        rom_memory[9891] = 3'b000;
        rom_memory[9892] = 3'b000;
        rom_memory[9893] = 3'b000;
        rom_memory[9894] = 3'b000;
        rom_memory[9895] = 3'b000;
        rom_memory[9896] = 3'b000;
        rom_memory[9897] = 3'b000;
        rom_memory[9898] = 3'b000;
        rom_memory[9899] = 3'b000;
        rom_memory[9900] = 3'b000;
        rom_memory[9901] = 3'b000;
        rom_memory[9902] = 3'b000;
        rom_memory[9903] = 3'b000;
        rom_memory[9904] = 3'b000;
        rom_memory[9905] = 3'b000;
        rom_memory[9906] = 3'b000;
        rom_memory[9907] = 3'b000;
        rom_memory[9908] = 3'b000;
        rom_memory[9909] = 3'b000;
        rom_memory[9910] = 3'b000;
        rom_memory[9911] = 3'b000;
        rom_memory[9912] = 3'b000;
        rom_memory[9913] = 3'b000;
        rom_memory[9914] = 3'b000;
        rom_memory[9915] = 3'b000;
        rom_memory[9916] = 3'b000;
        rom_memory[9917] = 3'b000;
        rom_memory[9918] = 3'b000;
        rom_memory[9919] = 3'b000;
        rom_memory[9920] = 3'b000;
        rom_memory[9921] = 3'b000;
        rom_memory[9922] = 3'b010;
        rom_memory[9923] = 3'b011;
        rom_memory[9924] = 3'b011;
        rom_memory[9925] = 3'b000;
        rom_memory[9926] = 3'b000;
        rom_memory[9927] = 3'b000;
        rom_memory[9928] = 3'b000;
        rom_memory[9929] = 3'b000;
        rom_memory[9930] = 3'b011;
        rom_memory[9931] = 3'b011;
        rom_memory[9932] = 3'b011;
        rom_memory[9933] = 3'b011;
        rom_memory[9934] = 3'b011;
        rom_memory[9935] = 3'b011;
        rom_memory[9936] = 3'b111;
        rom_memory[9937] = 3'b111;
        rom_memory[9938] = 3'b110;
        rom_memory[9939] = 3'b110;
        rom_memory[9940] = 3'b110;
        rom_memory[9941] = 3'b110;
        rom_memory[9942] = 3'b111;
        rom_memory[9943] = 3'b110;
        rom_memory[9944] = 3'b110;
        rom_memory[9945] = 3'b110;
        rom_memory[9946] = 3'b110;
        rom_memory[9947] = 3'b110;
        rom_memory[9948] = 3'b110;
        rom_memory[9949] = 3'b110;
        rom_memory[9950] = 3'b110;
        rom_memory[9951] = 3'b110;
        rom_memory[9952] = 3'b110;
        rom_memory[9953] = 3'b110;
        rom_memory[9954] = 3'b110;
        rom_memory[9955] = 3'b110;
        rom_memory[9956] = 3'b110;
        rom_memory[9957] = 3'b110;
        rom_memory[9958] = 3'b110;
        rom_memory[9959] = 3'b110;
        rom_memory[9960] = 3'b110;
        rom_memory[9961] = 3'b110;
        rom_memory[9962] = 3'b110;
        rom_memory[9963] = 3'b110;
        rom_memory[9964] = 3'b110;
        rom_memory[9965] = 3'b110;
        rom_memory[9966] = 3'b110;
        rom_memory[9967] = 3'b110;
        rom_memory[9968] = 3'b110;
        rom_memory[9969] = 3'b110;
        rom_memory[9970] = 3'b110;
        rom_memory[9971] = 3'b110;
        rom_memory[9972] = 3'b110;
        rom_memory[9973] = 3'b110;
        rom_memory[9974] = 3'b110;
        rom_memory[9975] = 3'b110;
        rom_memory[9976] = 3'b110;
        rom_memory[9977] = 3'b110;
        rom_memory[9978] = 3'b110;
        rom_memory[9979] = 3'b110;
        rom_memory[9980] = 3'b110;
        rom_memory[9981] = 3'b110;
        rom_memory[9982] = 3'b110;
        rom_memory[9983] = 3'b110;
        rom_memory[9984] = 3'b110;
        rom_memory[9985] = 3'b110;
        rom_memory[9986] = 3'b110;
        rom_memory[9987] = 3'b110;
        rom_memory[9988] = 3'b110;
        rom_memory[9989] = 3'b110;
        rom_memory[9990] = 3'b110;
        rom_memory[9991] = 3'b110;
        rom_memory[9992] = 3'b110;
        rom_memory[9993] = 3'b110;
        rom_memory[9994] = 3'b110;
        rom_memory[9995] = 3'b110;
        rom_memory[9996] = 3'b110;
        rom_memory[9997] = 3'b110;
        rom_memory[9998] = 3'b110;
        rom_memory[9999] = 3'b110;
        rom_memory[10000] = 3'b110;
        rom_memory[10001] = 3'b110;
        rom_memory[10002] = 3'b110;
        rom_memory[10003] = 3'b110;
        rom_memory[10004] = 3'b110;
        rom_memory[10005] = 3'b110;
        rom_memory[10006] = 3'b110;
        rom_memory[10007] = 3'b110;
        rom_memory[10008] = 3'b110;
        rom_memory[10009] = 3'b110;
        rom_memory[10010] = 3'b110;
        rom_memory[10011] = 3'b110;
        rom_memory[10012] = 3'b110;
        rom_memory[10013] = 3'b110;
        rom_memory[10014] = 3'b110;
        rom_memory[10015] = 3'b110;
        rom_memory[10016] = 3'b110;
        rom_memory[10017] = 3'b110;
        rom_memory[10018] = 3'b110;
        rom_memory[10019] = 3'b110;
        rom_memory[10020] = 3'b110;
        rom_memory[10021] = 3'b110;
        rom_memory[10022] = 3'b110;
        rom_memory[10023] = 3'b110;
        rom_memory[10024] = 3'b110;
        rom_memory[10025] = 3'b110;
        rom_memory[10026] = 3'b110;
        rom_memory[10027] = 3'b110;
        rom_memory[10028] = 3'b110;
        rom_memory[10029] = 3'b110;
        rom_memory[10030] = 3'b110;
        rom_memory[10031] = 3'b110;
        rom_memory[10032] = 3'b110;
        rom_memory[10033] = 3'b110;
        rom_memory[10034] = 3'b110;
        rom_memory[10035] = 3'b110;
        rom_memory[10036] = 3'b110;
        rom_memory[10037] = 3'b110;
        rom_memory[10038] = 3'b110;
        rom_memory[10039] = 3'b110;
        rom_memory[10040] = 3'b110;
        rom_memory[10041] = 3'b110;
        rom_memory[10042] = 3'b110;
        rom_memory[10043] = 3'b110;
        rom_memory[10044] = 3'b110;
        rom_memory[10045] = 3'b110;
        rom_memory[10046] = 3'b110;
        rom_memory[10047] = 3'b110;
        rom_memory[10048] = 3'b110;
        rom_memory[10049] = 3'b110;
        rom_memory[10050] = 3'b110;
        rom_memory[10051] = 3'b110;
        rom_memory[10052] = 3'b110;
        rom_memory[10053] = 3'b110;
        rom_memory[10054] = 3'b110;
        rom_memory[10055] = 3'b110;
        rom_memory[10056] = 3'b110;
        rom_memory[10057] = 3'b110;
        rom_memory[10058] = 3'b110;
        rom_memory[10059] = 3'b110;
        rom_memory[10060] = 3'b110;
        rom_memory[10061] = 3'b110;
        rom_memory[10062] = 3'b110;
        rom_memory[10063] = 3'b110;
        rom_memory[10064] = 3'b110;
        rom_memory[10065] = 3'b110;
        rom_memory[10066] = 3'b110;
        rom_memory[10067] = 3'b110;
        rom_memory[10068] = 3'b110;
        rom_memory[10069] = 3'b110;
        rom_memory[10070] = 3'b110;
        rom_memory[10071] = 3'b110;
        rom_memory[10072] = 3'b110;
        rom_memory[10073] = 3'b110;
        rom_memory[10074] = 3'b110;
        rom_memory[10075] = 3'b110;
        rom_memory[10076] = 3'b110;
        rom_memory[10077] = 3'b110;
        rom_memory[10078] = 3'b110;
        rom_memory[10079] = 3'b110;
        rom_memory[10080] = 3'b110;
        rom_memory[10081] = 3'b110;
        rom_memory[10082] = 3'b110;
        rom_memory[10083] = 3'b110;
        rom_memory[10084] = 3'b110;
        rom_memory[10085] = 3'b110;
        rom_memory[10086] = 3'b110;
        rom_memory[10087] = 3'b110;
        rom_memory[10088] = 3'b110;
        rom_memory[10089] = 3'b110;
        rom_memory[10090] = 3'b110;
        rom_memory[10091] = 3'b110;
        rom_memory[10092] = 3'b110;
        rom_memory[10093] = 3'b110;
        rom_memory[10094] = 3'b110;
        rom_memory[10095] = 3'b110;
        rom_memory[10096] = 3'b110;
        rom_memory[10097] = 3'b110;
        rom_memory[10098] = 3'b110;
        rom_memory[10099] = 3'b110;
        rom_memory[10100] = 3'b110;
        rom_memory[10101] = 3'b110;
        rom_memory[10102] = 3'b110;
        rom_memory[10103] = 3'b110;
        rom_memory[10104] = 3'b110;
        rom_memory[10105] = 3'b110;
        rom_memory[10106] = 3'b110;
        rom_memory[10107] = 3'b110;
        rom_memory[10108] = 3'b110;
        rom_memory[10109] = 3'b110;
        rom_memory[10110] = 3'b110;
        rom_memory[10111] = 3'b110;
        rom_memory[10112] = 3'b110;
        rom_memory[10113] = 3'b110;
        rom_memory[10114] = 3'b110;
        rom_memory[10115] = 3'b110;
        rom_memory[10116] = 3'b110;
        rom_memory[10117] = 3'b110;
        rom_memory[10118] = 3'b110;
        rom_memory[10119] = 3'b110;
        rom_memory[10120] = 3'b110;
        rom_memory[10121] = 3'b110;
        rom_memory[10122] = 3'b110;
        rom_memory[10123] = 3'b110;
        rom_memory[10124] = 3'b110;
        rom_memory[10125] = 3'b110;
        rom_memory[10126] = 3'b111;
        rom_memory[10127] = 3'b111;
        rom_memory[10128] = 3'b000;
        rom_memory[10129] = 3'b000;
        rom_memory[10130] = 3'b000;
        rom_memory[10131] = 3'b000;
        rom_memory[10132] = 3'b000;
        rom_memory[10133] = 3'b000;
        rom_memory[10134] = 3'b000;
        rom_memory[10135] = 3'b000;
        rom_memory[10136] = 3'b000;
        rom_memory[10137] = 3'b000;
        rom_memory[10138] = 3'b000;
        rom_memory[10139] = 3'b000;
        rom_memory[10140] = 3'b000;
        rom_memory[10141] = 3'b000;
        rom_memory[10142] = 3'b000;
        rom_memory[10143] = 3'b000;
        rom_memory[10144] = 3'b000;
        rom_memory[10145] = 3'b000;
        rom_memory[10146] = 3'b000;
        rom_memory[10147] = 3'b000;
        rom_memory[10148] = 3'b000;
        rom_memory[10149] = 3'b000;
        rom_memory[10150] = 3'b000;
        rom_memory[10151] = 3'b000;
        rom_memory[10152] = 3'b000;
        rom_memory[10153] = 3'b000;
        rom_memory[10154] = 3'b000;
        rom_memory[10155] = 3'b000;
        rom_memory[10156] = 3'b000;
        rom_memory[10157] = 3'b000;
        rom_memory[10158] = 3'b000;
        rom_memory[10159] = 3'b000;
        rom_memory[10160] = 3'b000;
        rom_memory[10161] = 3'b000;
        rom_memory[10162] = 3'b000;
        rom_memory[10163] = 3'b000;
        rom_memory[10164] = 3'b011;
        rom_memory[10165] = 3'b000;
        rom_memory[10166] = 3'b000;
        rom_memory[10167] = 3'b010;
        rom_memory[10168] = 3'b011;
        rom_memory[10169] = 3'b011;
        rom_memory[10170] = 3'b011;
        rom_memory[10171] = 3'b011;
        rom_memory[10172] = 3'b011;
        rom_memory[10173] = 3'b011;
        rom_memory[10174] = 3'b011;
        rom_memory[10175] = 3'b011;
        rom_memory[10176] = 3'b011;
        rom_memory[10177] = 3'b111;
        rom_memory[10178] = 3'b111;
        rom_memory[10179] = 3'b110;
        rom_memory[10180] = 3'b110;
        rom_memory[10181] = 3'b110;
        rom_memory[10182] = 3'b110;
        rom_memory[10183] = 3'b110;
        rom_memory[10184] = 3'b110;
        rom_memory[10185] = 3'b110;
        rom_memory[10186] = 3'b110;
        rom_memory[10187] = 3'b110;
        rom_memory[10188] = 3'b110;
        rom_memory[10189] = 3'b110;
        rom_memory[10190] = 3'b110;
        rom_memory[10191] = 3'b110;
        rom_memory[10192] = 3'b110;
        rom_memory[10193] = 3'b110;
        rom_memory[10194] = 3'b110;
        rom_memory[10195] = 3'b110;
        rom_memory[10196] = 3'b110;
        rom_memory[10197] = 3'b110;
        rom_memory[10198] = 3'b110;
        rom_memory[10199] = 3'b110;
        rom_memory[10200] = 3'b110;
        rom_memory[10201] = 3'b110;
        rom_memory[10202] = 3'b110;
        rom_memory[10203] = 3'b110;
        rom_memory[10204] = 3'b110;
        rom_memory[10205] = 3'b110;
        rom_memory[10206] = 3'b110;
        rom_memory[10207] = 3'b110;
        rom_memory[10208] = 3'b110;
        rom_memory[10209] = 3'b110;
        rom_memory[10210] = 3'b110;
        rom_memory[10211] = 3'b110;
        rom_memory[10212] = 3'b110;
        rom_memory[10213] = 3'b110;
        rom_memory[10214] = 3'b110;
        rom_memory[10215] = 3'b110;
        rom_memory[10216] = 3'b110;
        rom_memory[10217] = 3'b110;
        rom_memory[10218] = 3'b110;
        rom_memory[10219] = 3'b110;
        rom_memory[10220] = 3'b110;
        rom_memory[10221] = 3'b110;
        rom_memory[10222] = 3'b110;
        rom_memory[10223] = 3'b110;
        rom_memory[10224] = 3'b110;
        rom_memory[10225] = 3'b110;
        rom_memory[10226] = 3'b110;
        rom_memory[10227] = 3'b110;
        rom_memory[10228] = 3'b110;
        rom_memory[10229] = 3'b110;
        rom_memory[10230] = 3'b110;
        rom_memory[10231] = 3'b110;
        rom_memory[10232] = 3'b110;
        rom_memory[10233] = 3'b110;
        rom_memory[10234] = 3'b110;
        rom_memory[10235] = 3'b110;
        rom_memory[10236] = 3'b110;
        rom_memory[10237] = 3'b110;
        rom_memory[10238] = 3'b110;
        rom_memory[10239] = 3'b110;
        rom_memory[10240] = 3'b110;
        rom_memory[10241] = 3'b110;
        rom_memory[10242] = 3'b110;
        rom_memory[10243] = 3'b110;
        rom_memory[10244] = 3'b110;
        rom_memory[10245] = 3'b110;
        rom_memory[10246] = 3'b110;
        rom_memory[10247] = 3'b110;
        rom_memory[10248] = 3'b110;
        rom_memory[10249] = 3'b110;
        rom_memory[10250] = 3'b110;
        rom_memory[10251] = 3'b110;
        rom_memory[10252] = 3'b110;
        rom_memory[10253] = 3'b110;
        rom_memory[10254] = 3'b110;
        rom_memory[10255] = 3'b110;
        rom_memory[10256] = 3'b110;
        rom_memory[10257] = 3'b110;
        rom_memory[10258] = 3'b110;
        rom_memory[10259] = 3'b110;
        rom_memory[10260] = 3'b110;
        rom_memory[10261] = 3'b110;
        rom_memory[10262] = 3'b110;
        rom_memory[10263] = 3'b110;
        rom_memory[10264] = 3'b110;
        rom_memory[10265] = 3'b110;
        rom_memory[10266] = 3'b110;
        rom_memory[10267] = 3'b110;
        rom_memory[10268] = 3'b110;
        rom_memory[10269] = 3'b110;
        rom_memory[10270] = 3'b110;
        rom_memory[10271] = 3'b110;
        rom_memory[10272] = 3'b110;
        rom_memory[10273] = 3'b110;
        rom_memory[10274] = 3'b110;
        rom_memory[10275] = 3'b110;
        rom_memory[10276] = 3'b110;
        rom_memory[10277] = 3'b110;
        rom_memory[10278] = 3'b110;
        rom_memory[10279] = 3'b110;
        rom_memory[10280] = 3'b110;
        rom_memory[10281] = 3'b110;
        rom_memory[10282] = 3'b110;
        rom_memory[10283] = 3'b110;
        rom_memory[10284] = 3'b110;
        rom_memory[10285] = 3'b110;
        rom_memory[10286] = 3'b110;
        rom_memory[10287] = 3'b110;
        rom_memory[10288] = 3'b110;
        rom_memory[10289] = 3'b110;
        rom_memory[10290] = 3'b110;
        rom_memory[10291] = 3'b110;
        rom_memory[10292] = 3'b110;
        rom_memory[10293] = 3'b110;
        rom_memory[10294] = 3'b110;
        rom_memory[10295] = 3'b110;
        rom_memory[10296] = 3'b110;
        rom_memory[10297] = 3'b110;
        rom_memory[10298] = 3'b110;
        rom_memory[10299] = 3'b110;
        rom_memory[10300] = 3'b110;
        rom_memory[10301] = 3'b110;
        rom_memory[10302] = 3'b110;
        rom_memory[10303] = 3'b110;
        rom_memory[10304] = 3'b110;
        rom_memory[10305] = 3'b110;
        rom_memory[10306] = 3'b110;
        rom_memory[10307] = 3'b110;
        rom_memory[10308] = 3'b110;
        rom_memory[10309] = 3'b110;
        rom_memory[10310] = 3'b110;
        rom_memory[10311] = 3'b110;
        rom_memory[10312] = 3'b110;
        rom_memory[10313] = 3'b110;
        rom_memory[10314] = 3'b110;
        rom_memory[10315] = 3'b110;
        rom_memory[10316] = 3'b110;
        rom_memory[10317] = 3'b110;
        rom_memory[10318] = 3'b110;
        rom_memory[10319] = 3'b110;
        rom_memory[10320] = 3'b110;
        rom_memory[10321] = 3'b110;
        rom_memory[10322] = 3'b110;
        rom_memory[10323] = 3'b110;
        rom_memory[10324] = 3'b110;
        rom_memory[10325] = 3'b110;
        rom_memory[10326] = 3'b110;
        rom_memory[10327] = 3'b110;
        rom_memory[10328] = 3'b110;
        rom_memory[10329] = 3'b110;
        rom_memory[10330] = 3'b110;
        rom_memory[10331] = 3'b110;
        rom_memory[10332] = 3'b110;
        rom_memory[10333] = 3'b110;
        rom_memory[10334] = 3'b110;
        rom_memory[10335] = 3'b110;
        rom_memory[10336] = 3'b110;
        rom_memory[10337] = 3'b110;
        rom_memory[10338] = 3'b110;
        rom_memory[10339] = 3'b110;
        rom_memory[10340] = 3'b110;
        rom_memory[10341] = 3'b110;
        rom_memory[10342] = 3'b110;
        rom_memory[10343] = 3'b110;
        rom_memory[10344] = 3'b110;
        rom_memory[10345] = 3'b110;
        rom_memory[10346] = 3'b110;
        rom_memory[10347] = 3'b110;
        rom_memory[10348] = 3'b110;
        rom_memory[10349] = 3'b110;
        rom_memory[10350] = 3'b110;
        rom_memory[10351] = 3'b110;
        rom_memory[10352] = 3'b110;
        rom_memory[10353] = 3'b110;
        rom_memory[10354] = 3'b110;
        rom_memory[10355] = 3'b110;
        rom_memory[10356] = 3'b110;
        rom_memory[10357] = 3'b110;
        rom_memory[10358] = 3'b110;
        rom_memory[10359] = 3'b110;
        rom_memory[10360] = 3'b110;
        rom_memory[10361] = 3'b110;
        rom_memory[10362] = 3'b110;
        rom_memory[10363] = 3'b110;
        rom_memory[10364] = 3'b110;
        rom_memory[10365] = 3'b111;
        rom_memory[10366] = 3'b111;
        rom_memory[10367] = 3'b110;
        rom_memory[10368] = 3'b000;
        rom_memory[10369] = 3'b000;
        rom_memory[10370] = 3'b000;
        rom_memory[10371] = 3'b000;
        rom_memory[10372] = 3'b000;
        rom_memory[10373] = 3'b000;
        rom_memory[10374] = 3'b000;
        rom_memory[10375] = 3'b000;
        rom_memory[10376] = 3'b000;
        rom_memory[10377] = 3'b000;
        rom_memory[10378] = 3'b000;
        rom_memory[10379] = 3'b000;
        rom_memory[10380] = 3'b000;
        rom_memory[10381] = 3'b000;
        rom_memory[10382] = 3'b000;
        rom_memory[10383] = 3'b000;
        rom_memory[10384] = 3'b000;
        rom_memory[10385] = 3'b000;
        rom_memory[10386] = 3'b000;
        rom_memory[10387] = 3'b000;
        rom_memory[10388] = 3'b000;
        rom_memory[10389] = 3'b000;
        rom_memory[10390] = 3'b000;
        rom_memory[10391] = 3'b000;
        rom_memory[10392] = 3'b000;
        rom_memory[10393] = 3'b000;
        rom_memory[10394] = 3'b000;
        rom_memory[10395] = 3'b000;
        rom_memory[10396] = 3'b000;
        rom_memory[10397] = 3'b000;
        rom_memory[10398] = 3'b000;
        rom_memory[10399] = 3'b000;
        rom_memory[10400] = 3'b000;
        rom_memory[10401] = 3'b000;
        rom_memory[10402] = 3'b000;
        rom_memory[10403] = 3'b000;
        rom_memory[10404] = 3'b000;
        rom_memory[10405] = 3'b011;
        rom_memory[10406] = 3'b011;
        rom_memory[10407] = 3'b011;
        rom_memory[10408] = 3'b011;
        rom_memory[10409] = 3'b011;
        rom_memory[10410] = 3'b011;
        rom_memory[10411] = 3'b000;
        rom_memory[10412] = 3'b011;
        rom_memory[10413] = 3'b011;
        rom_memory[10414] = 3'b011;
        rom_memory[10415] = 3'b011;
        rom_memory[10416] = 3'b011;
        rom_memory[10417] = 3'b001;
        rom_memory[10418] = 3'b111;
        rom_memory[10419] = 3'b110;
        rom_memory[10420] = 3'b110;
        rom_memory[10421] = 3'b110;
        rom_memory[10422] = 3'b110;
        rom_memory[10423] = 3'b110;
        rom_memory[10424] = 3'b110;
        rom_memory[10425] = 3'b110;
        rom_memory[10426] = 3'b110;
        rom_memory[10427] = 3'b110;
        rom_memory[10428] = 3'b110;
        rom_memory[10429] = 3'b110;
        rom_memory[10430] = 3'b110;
        rom_memory[10431] = 3'b110;
        rom_memory[10432] = 3'b110;
        rom_memory[10433] = 3'b110;
        rom_memory[10434] = 3'b110;
        rom_memory[10435] = 3'b110;
        rom_memory[10436] = 3'b110;
        rom_memory[10437] = 3'b110;
        rom_memory[10438] = 3'b110;
        rom_memory[10439] = 3'b110;
        rom_memory[10440] = 3'b110;
        rom_memory[10441] = 3'b110;
        rom_memory[10442] = 3'b110;
        rom_memory[10443] = 3'b110;
        rom_memory[10444] = 3'b110;
        rom_memory[10445] = 3'b110;
        rom_memory[10446] = 3'b110;
        rom_memory[10447] = 3'b110;
        rom_memory[10448] = 3'b110;
        rom_memory[10449] = 3'b110;
        rom_memory[10450] = 3'b110;
        rom_memory[10451] = 3'b110;
        rom_memory[10452] = 3'b110;
        rom_memory[10453] = 3'b110;
        rom_memory[10454] = 3'b110;
        rom_memory[10455] = 3'b110;
        rom_memory[10456] = 3'b110;
        rom_memory[10457] = 3'b110;
        rom_memory[10458] = 3'b110;
        rom_memory[10459] = 3'b110;
        rom_memory[10460] = 3'b110;
        rom_memory[10461] = 3'b110;
        rom_memory[10462] = 3'b110;
        rom_memory[10463] = 3'b110;
        rom_memory[10464] = 3'b110;
        rom_memory[10465] = 3'b110;
        rom_memory[10466] = 3'b110;
        rom_memory[10467] = 3'b110;
        rom_memory[10468] = 3'b110;
        rom_memory[10469] = 3'b110;
        rom_memory[10470] = 3'b110;
        rom_memory[10471] = 3'b110;
        rom_memory[10472] = 3'b110;
        rom_memory[10473] = 3'b110;
        rom_memory[10474] = 3'b110;
        rom_memory[10475] = 3'b110;
        rom_memory[10476] = 3'b110;
        rom_memory[10477] = 3'b110;
        rom_memory[10478] = 3'b110;
        rom_memory[10479] = 3'b110;
        rom_memory[10480] = 3'b110;
        rom_memory[10481] = 3'b110;
        rom_memory[10482] = 3'b110;
        rom_memory[10483] = 3'b110;
        rom_memory[10484] = 3'b110;
        rom_memory[10485] = 3'b110;
        rom_memory[10486] = 3'b110;
        rom_memory[10487] = 3'b110;
        rom_memory[10488] = 3'b110;
        rom_memory[10489] = 3'b110;
        rom_memory[10490] = 3'b110;
        rom_memory[10491] = 3'b110;
        rom_memory[10492] = 3'b110;
        rom_memory[10493] = 3'b110;
        rom_memory[10494] = 3'b110;
        rom_memory[10495] = 3'b110;
        rom_memory[10496] = 3'b110;
        rom_memory[10497] = 3'b110;
        rom_memory[10498] = 3'b110;
        rom_memory[10499] = 3'b110;
        rom_memory[10500] = 3'b110;
        rom_memory[10501] = 3'b110;
        rom_memory[10502] = 3'b110;
        rom_memory[10503] = 3'b110;
        rom_memory[10504] = 3'b110;
        rom_memory[10505] = 3'b110;
        rom_memory[10506] = 3'b110;
        rom_memory[10507] = 3'b110;
        rom_memory[10508] = 3'b110;
        rom_memory[10509] = 3'b110;
        rom_memory[10510] = 3'b110;
        rom_memory[10511] = 3'b110;
        rom_memory[10512] = 3'b110;
        rom_memory[10513] = 3'b110;
        rom_memory[10514] = 3'b110;
        rom_memory[10515] = 3'b110;
        rom_memory[10516] = 3'b110;
        rom_memory[10517] = 3'b110;
        rom_memory[10518] = 3'b110;
        rom_memory[10519] = 3'b110;
        rom_memory[10520] = 3'b110;
        rom_memory[10521] = 3'b110;
        rom_memory[10522] = 3'b110;
        rom_memory[10523] = 3'b110;
        rom_memory[10524] = 3'b110;
        rom_memory[10525] = 3'b110;
        rom_memory[10526] = 3'b110;
        rom_memory[10527] = 3'b110;
        rom_memory[10528] = 3'b110;
        rom_memory[10529] = 3'b110;
        rom_memory[10530] = 3'b110;
        rom_memory[10531] = 3'b110;
        rom_memory[10532] = 3'b110;
        rom_memory[10533] = 3'b110;
        rom_memory[10534] = 3'b110;
        rom_memory[10535] = 3'b110;
        rom_memory[10536] = 3'b110;
        rom_memory[10537] = 3'b110;
        rom_memory[10538] = 3'b110;
        rom_memory[10539] = 3'b110;
        rom_memory[10540] = 3'b110;
        rom_memory[10541] = 3'b110;
        rom_memory[10542] = 3'b110;
        rom_memory[10543] = 3'b110;
        rom_memory[10544] = 3'b110;
        rom_memory[10545] = 3'b110;
        rom_memory[10546] = 3'b110;
        rom_memory[10547] = 3'b110;
        rom_memory[10548] = 3'b110;
        rom_memory[10549] = 3'b110;
        rom_memory[10550] = 3'b110;
        rom_memory[10551] = 3'b110;
        rom_memory[10552] = 3'b110;
        rom_memory[10553] = 3'b110;
        rom_memory[10554] = 3'b110;
        rom_memory[10555] = 3'b110;
        rom_memory[10556] = 3'b110;
        rom_memory[10557] = 3'b110;
        rom_memory[10558] = 3'b110;
        rom_memory[10559] = 3'b110;
        rom_memory[10560] = 3'b110;
        rom_memory[10561] = 3'b110;
        rom_memory[10562] = 3'b110;
        rom_memory[10563] = 3'b110;
        rom_memory[10564] = 3'b110;
        rom_memory[10565] = 3'b110;
        rom_memory[10566] = 3'b110;
        rom_memory[10567] = 3'b110;
        rom_memory[10568] = 3'b110;
        rom_memory[10569] = 3'b110;
        rom_memory[10570] = 3'b110;
        rom_memory[10571] = 3'b110;
        rom_memory[10572] = 3'b110;
        rom_memory[10573] = 3'b110;
        rom_memory[10574] = 3'b110;
        rom_memory[10575] = 3'b110;
        rom_memory[10576] = 3'b110;
        rom_memory[10577] = 3'b110;
        rom_memory[10578] = 3'b110;
        rom_memory[10579] = 3'b110;
        rom_memory[10580] = 3'b110;
        rom_memory[10581] = 3'b110;
        rom_memory[10582] = 3'b110;
        rom_memory[10583] = 3'b110;
        rom_memory[10584] = 3'b110;
        rom_memory[10585] = 3'b110;
        rom_memory[10586] = 3'b110;
        rom_memory[10587] = 3'b110;
        rom_memory[10588] = 3'b110;
        rom_memory[10589] = 3'b110;
        rom_memory[10590] = 3'b110;
        rom_memory[10591] = 3'b110;
        rom_memory[10592] = 3'b110;
        rom_memory[10593] = 3'b110;
        rom_memory[10594] = 3'b110;
        rom_memory[10595] = 3'b110;
        rom_memory[10596] = 3'b110;
        rom_memory[10597] = 3'b110;
        rom_memory[10598] = 3'b110;
        rom_memory[10599] = 3'b110;
        rom_memory[10600] = 3'b110;
        rom_memory[10601] = 3'b110;
        rom_memory[10602] = 3'b110;
        rom_memory[10603] = 3'b110;
        rom_memory[10604] = 3'b110;
        rom_memory[10605] = 3'b111;
        rom_memory[10606] = 3'b111;
        rom_memory[10607] = 3'b110;
        rom_memory[10608] = 3'b000;
        rom_memory[10609] = 3'b000;
        rom_memory[10610] = 3'b000;
        rom_memory[10611] = 3'b000;
        rom_memory[10612] = 3'b000;
        rom_memory[10613] = 3'b000;
        rom_memory[10614] = 3'b000;
        rom_memory[10615] = 3'b000;
        rom_memory[10616] = 3'b000;
        rom_memory[10617] = 3'b000;
        rom_memory[10618] = 3'b000;
        rom_memory[10619] = 3'b000;
        rom_memory[10620] = 3'b000;
        rom_memory[10621] = 3'b000;
        rom_memory[10622] = 3'b000;
        rom_memory[10623] = 3'b000;
        rom_memory[10624] = 3'b000;
        rom_memory[10625] = 3'b000;
        rom_memory[10626] = 3'b000;
        rom_memory[10627] = 3'b000;
        rom_memory[10628] = 3'b000;
        rom_memory[10629] = 3'b000;
        rom_memory[10630] = 3'b000;
        rom_memory[10631] = 3'b000;
        rom_memory[10632] = 3'b000;
        rom_memory[10633] = 3'b000;
        rom_memory[10634] = 3'b000;
        rom_memory[10635] = 3'b000;
        rom_memory[10636] = 3'b000;
        rom_memory[10637] = 3'b000;
        rom_memory[10638] = 3'b000;
        rom_memory[10639] = 3'b000;
        rom_memory[10640] = 3'b000;
        rom_memory[10641] = 3'b000;
        rom_memory[10642] = 3'b000;
        rom_memory[10643] = 3'b000;
        rom_memory[10644] = 3'b000;
        rom_memory[10645] = 3'b011;
        rom_memory[10646] = 3'b011;
        rom_memory[10647] = 3'b011;
        rom_memory[10648] = 3'b011;
        rom_memory[10649] = 3'b000;
        rom_memory[10650] = 3'b000;
        rom_memory[10651] = 3'b011;
        rom_memory[10652] = 3'b011;
        rom_memory[10653] = 3'b011;
        rom_memory[10654] = 3'b011;
        rom_memory[10655] = 3'b011;
        rom_memory[10656] = 3'b011;
        rom_memory[10657] = 3'b011;
        rom_memory[10658] = 3'b111;
        rom_memory[10659] = 3'b111;
        rom_memory[10660] = 3'b110;
        rom_memory[10661] = 3'b110;
        rom_memory[10662] = 3'b110;
        rom_memory[10663] = 3'b110;
        rom_memory[10664] = 3'b110;
        rom_memory[10665] = 3'b110;
        rom_memory[10666] = 3'b110;
        rom_memory[10667] = 3'b110;
        rom_memory[10668] = 3'b110;
        rom_memory[10669] = 3'b110;
        rom_memory[10670] = 3'b110;
        rom_memory[10671] = 3'b110;
        rom_memory[10672] = 3'b110;
        rom_memory[10673] = 3'b110;
        rom_memory[10674] = 3'b110;
        rom_memory[10675] = 3'b110;
        rom_memory[10676] = 3'b110;
        rom_memory[10677] = 3'b110;
        rom_memory[10678] = 3'b110;
        rom_memory[10679] = 3'b110;
        rom_memory[10680] = 3'b110;
        rom_memory[10681] = 3'b110;
        rom_memory[10682] = 3'b110;
        rom_memory[10683] = 3'b110;
        rom_memory[10684] = 3'b110;
        rom_memory[10685] = 3'b110;
        rom_memory[10686] = 3'b110;
        rom_memory[10687] = 3'b110;
        rom_memory[10688] = 3'b110;
        rom_memory[10689] = 3'b110;
        rom_memory[10690] = 3'b110;
        rom_memory[10691] = 3'b110;
        rom_memory[10692] = 3'b110;
        rom_memory[10693] = 3'b110;
        rom_memory[10694] = 3'b110;
        rom_memory[10695] = 3'b110;
        rom_memory[10696] = 3'b110;
        rom_memory[10697] = 3'b110;
        rom_memory[10698] = 3'b110;
        rom_memory[10699] = 3'b110;
        rom_memory[10700] = 3'b110;
        rom_memory[10701] = 3'b110;
        rom_memory[10702] = 3'b110;
        rom_memory[10703] = 3'b110;
        rom_memory[10704] = 3'b110;
        rom_memory[10705] = 3'b110;
        rom_memory[10706] = 3'b110;
        rom_memory[10707] = 3'b110;
        rom_memory[10708] = 3'b110;
        rom_memory[10709] = 3'b110;
        rom_memory[10710] = 3'b110;
        rom_memory[10711] = 3'b110;
        rom_memory[10712] = 3'b110;
        rom_memory[10713] = 3'b110;
        rom_memory[10714] = 3'b110;
        rom_memory[10715] = 3'b110;
        rom_memory[10716] = 3'b110;
        rom_memory[10717] = 3'b110;
        rom_memory[10718] = 3'b110;
        rom_memory[10719] = 3'b110;
        rom_memory[10720] = 3'b110;
        rom_memory[10721] = 3'b110;
        rom_memory[10722] = 3'b110;
        rom_memory[10723] = 3'b110;
        rom_memory[10724] = 3'b110;
        rom_memory[10725] = 3'b110;
        rom_memory[10726] = 3'b110;
        rom_memory[10727] = 3'b110;
        rom_memory[10728] = 3'b110;
        rom_memory[10729] = 3'b110;
        rom_memory[10730] = 3'b110;
        rom_memory[10731] = 3'b110;
        rom_memory[10732] = 3'b110;
        rom_memory[10733] = 3'b110;
        rom_memory[10734] = 3'b110;
        rom_memory[10735] = 3'b110;
        rom_memory[10736] = 3'b110;
        rom_memory[10737] = 3'b110;
        rom_memory[10738] = 3'b110;
        rom_memory[10739] = 3'b110;
        rom_memory[10740] = 3'b110;
        rom_memory[10741] = 3'b110;
        rom_memory[10742] = 3'b110;
        rom_memory[10743] = 3'b110;
        rom_memory[10744] = 3'b110;
        rom_memory[10745] = 3'b110;
        rom_memory[10746] = 3'b110;
        rom_memory[10747] = 3'b110;
        rom_memory[10748] = 3'b110;
        rom_memory[10749] = 3'b110;
        rom_memory[10750] = 3'b110;
        rom_memory[10751] = 3'b110;
        rom_memory[10752] = 3'b110;
        rom_memory[10753] = 3'b110;
        rom_memory[10754] = 3'b110;
        rom_memory[10755] = 3'b110;
        rom_memory[10756] = 3'b110;
        rom_memory[10757] = 3'b110;
        rom_memory[10758] = 3'b110;
        rom_memory[10759] = 3'b110;
        rom_memory[10760] = 3'b110;
        rom_memory[10761] = 3'b110;
        rom_memory[10762] = 3'b110;
        rom_memory[10763] = 3'b110;
        rom_memory[10764] = 3'b110;
        rom_memory[10765] = 3'b110;
        rom_memory[10766] = 3'b110;
        rom_memory[10767] = 3'b110;
        rom_memory[10768] = 3'b110;
        rom_memory[10769] = 3'b110;
        rom_memory[10770] = 3'b110;
        rom_memory[10771] = 3'b110;
        rom_memory[10772] = 3'b110;
        rom_memory[10773] = 3'b110;
        rom_memory[10774] = 3'b110;
        rom_memory[10775] = 3'b110;
        rom_memory[10776] = 3'b110;
        rom_memory[10777] = 3'b110;
        rom_memory[10778] = 3'b110;
        rom_memory[10779] = 3'b110;
        rom_memory[10780] = 3'b110;
        rom_memory[10781] = 3'b110;
        rom_memory[10782] = 3'b110;
        rom_memory[10783] = 3'b110;
        rom_memory[10784] = 3'b110;
        rom_memory[10785] = 3'b110;
        rom_memory[10786] = 3'b110;
        rom_memory[10787] = 3'b110;
        rom_memory[10788] = 3'b110;
        rom_memory[10789] = 3'b110;
        rom_memory[10790] = 3'b110;
        rom_memory[10791] = 3'b110;
        rom_memory[10792] = 3'b110;
        rom_memory[10793] = 3'b110;
        rom_memory[10794] = 3'b110;
        rom_memory[10795] = 3'b110;
        rom_memory[10796] = 3'b110;
        rom_memory[10797] = 3'b110;
        rom_memory[10798] = 3'b110;
        rom_memory[10799] = 3'b110;
        rom_memory[10800] = 3'b110;
        rom_memory[10801] = 3'b110;
        rom_memory[10802] = 3'b110;
        rom_memory[10803] = 3'b110;
        rom_memory[10804] = 3'b110;
        rom_memory[10805] = 3'b110;
        rom_memory[10806] = 3'b110;
        rom_memory[10807] = 3'b110;
        rom_memory[10808] = 3'b110;
        rom_memory[10809] = 3'b110;
        rom_memory[10810] = 3'b110;
        rom_memory[10811] = 3'b110;
        rom_memory[10812] = 3'b110;
        rom_memory[10813] = 3'b110;
        rom_memory[10814] = 3'b110;
        rom_memory[10815] = 3'b110;
        rom_memory[10816] = 3'b110;
        rom_memory[10817] = 3'b110;
        rom_memory[10818] = 3'b110;
        rom_memory[10819] = 3'b110;
        rom_memory[10820] = 3'b110;
        rom_memory[10821] = 3'b110;
        rom_memory[10822] = 3'b110;
        rom_memory[10823] = 3'b110;
        rom_memory[10824] = 3'b110;
        rom_memory[10825] = 3'b110;
        rom_memory[10826] = 3'b110;
        rom_memory[10827] = 3'b110;
        rom_memory[10828] = 3'b110;
        rom_memory[10829] = 3'b110;
        rom_memory[10830] = 3'b110;
        rom_memory[10831] = 3'b110;
        rom_memory[10832] = 3'b110;
        rom_memory[10833] = 3'b110;
        rom_memory[10834] = 3'b110;
        rom_memory[10835] = 3'b110;
        rom_memory[10836] = 3'b110;
        rom_memory[10837] = 3'b110;
        rom_memory[10838] = 3'b110;
        rom_memory[10839] = 3'b110;
        rom_memory[10840] = 3'b110;
        rom_memory[10841] = 3'b110;
        rom_memory[10842] = 3'b110;
        rom_memory[10843] = 3'b110;
        rom_memory[10844] = 3'b110;
        rom_memory[10845] = 3'b111;
        rom_memory[10846] = 3'b111;
        rom_memory[10847] = 3'b111;
        rom_memory[10848] = 3'b000;
        rom_memory[10849] = 3'b000;
        rom_memory[10850] = 3'b000;
        rom_memory[10851] = 3'b000;
        rom_memory[10852] = 3'b000;
        rom_memory[10853] = 3'b000;
        rom_memory[10854] = 3'b000;
        rom_memory[10855] = 3'b000;
        rom_memory[10856] = 3'b000;
        rom_memory[10857] = 3'b000;
        rom_memory[10858] = 3'b000;
        rom_memory[10859] = 3'b000;
        rom_memory[10860] = 3'b000;
        rom_memory[10861] = 3'b000;
        rom_memory[10862] = 3'b000;
        rom_memory[10863] = 3'b000;
        rom_memory[10864] = 3'b000;
        rom_memory[10865] = 3'b000;
        rom_memory[10866] = 3'b000;
        rom_memory[10867] = 3'b000;
        rom_memory[10868] = 3'b000;
        rom_memory[10869] = 3'b000;
        rom_memory[10870] = 3'b000;
        rom_memory[10871] = 3'b000;
        rom_memory[10872] = 3'b000;
        rom_memory[10873] = 3'b000;
        rom_memory[10874] = 3'b000;
        rom_memory[10875] = 3'b000;
        rom_memory[10876] = 3'b000;
        rom_memory[10877] = 3'b000;
        rom_memory[10878] = 3'b000;
        rom_memory[10879] = 3'b000;
        rom_memory[10880] = 3'b000;
        rom_memory[10881] = 3'b000;
        rom_memory[10882] = 3'b000;
        rom_memory[10883] = 3'b000;
        rom_memory[10884] = 3'b000;
        rom_memory[10885] = 3'b000;
        rom_memory[10886] = 3'b011;
        rom_memory[10887] = 3'b011;
        rom_memory[10888] = 3'b011;
        rom_memory[10889] = 3'b011;
        rom_memory[10890] = 3'b011;
        rom_memory[10891] = 3'b011;
        rom_memory[10892] = 3'b001;
        rom_memory[10893] = 3'b011;
        rom_memory[10894] = 3'b011;
        rom_memory[10895] = 3'b011;
        rom_memory[10896] = 3'b011;
        rom_memory[10897] = 3'b111;
        rom_memory[10898] = 3'b111;
        rom_memory[10899] = 3'b111;
        rom_memory[10900] = 3'b111;
        rom_memory[10901] = 3'b110;
        rom_memory[10902] = 3'b110;
        rom_memory[10903] = 3'b110;
        rom_memory[10904] = 3'b110;
        rom_memory[10905] = 3'b110;
        rom_memory[10906] = 3'b110;
        rom_memory[10907] = 3'b110;
        rom_memory[10908] = 3'b110;
        rom_memory[10909] = 3'b110;
        rom_memory[10910] = 3'b110;
        rom_memory[10911] = 3'b110;
        rom_memory[10912] = 3'b110;
        rom_memory[10913] = 3'b110;
        rom_memory[10914] = 3'b110;
        rom_memory[10915] = 3'b110;
        rom_memory[10916] = 3'b110;
        rom_memory[10917] = 3'b110;
        rom_memory[10918] = 3'b110;
        rom_memory[10919] = 3'b110;
        rom_memory[10920] = 3'b110;
        rom_memory[10921] = 3'b110;
        rom_memory[10922] = 3'b110;
        rom_memory[10923] = 3'b110;
        rom_memory[10924] = 3'b110;
        rom_memory[10925] = 3'b110;
        rom_memory[10926] = 3'b110;
        rom_memory[10927] = 3'b110;
        rom_memory[10928] = 3'b110;
        rom_memory[10929] = 3'b110;
        rom_memory[10930] = 3'b110;
        rom_memory[10931] = 3'b110;
        rom_memory[10932] = 3'b110;
        rom_memory[10933] = 3'b110;
        rom_memory[10934] = 3'b110;
        rom_memory[10935] = 3'b110;
        rom_memory[10936] = 3'b110;
        rom_memory[10937] = 3'b110;
        rom_memory[10938] = 3'b110;
        rom_memory[10939] = 3'b110;
        rom_memory[10940] = 3'b110;
        rom_memory[10941] = 3'b110;
        rom_memory[10942] = 3'b110;
        rom_memory[10943] = 3'b110;
        rom_memory[10944] = 3'b110;
        rom_memory[10945] = 3'b110;
        rom_memory[10946] = 3'b110;
        rom_memory[10947] = 3'b110;
        rom_memory[10948] = 3'b110;
        rom_memory[10949] = 3'b110;
        rom_memory[10950] = 3'b110;
        rom_memory[10951] = 3'b110;
        rom_memory[10952] = 3'b110;
        rom_memory[10953] = 3'b110;
        rom_memory[10954] = 3'b110;
        rom_memory[10955] = 3'b110;
        rom_memory[10956] = 3'b110;
        rom_memory[10957] = 3'b110;
        rom_memory[10958] = 3'b110;
        rom_memory[10959] = 3'b110;
        rom_memory[10960] = 3'b110;
        rom_memory[10961] = 3'b110;
        rom_memory[10962] = 3'b110;
        rom_memory[10963] = 3'b110;
        rom_memory[10964] = 3'b110;
        rom_memory[10965] = 3'b110;
        rom_memory[10966] = 3'b110;
        rom_memory[10967] = 3'b110;
        rom_memory[10968] = 3'b110;
        rom_memory[10969] = 3'b110;
        rom_memory[10970] = 3'b110;
        rom_memory[10971] = 3'b110;
        rom_memory[10972] = 3'b110;
        rom_memory[10973] = 3'b110;
        rom_memory[10974] = 3'b110;
        rom_memory[10975] = 3'b110;
        rom_memory[10976] = 3'b110;
        rom_memory[10977] = 3'b110;
        rom_memory[10978] = 3'b110;
        rom_memory[10979] = 3'b110;
        rom_memory[10980] = 3'b110;
        rom_memory[10981] = 3'b110;
        rom_memory[10982] = 3'b110;
        rom_memory[10983] = 3'b110;
        rom_memory[10984] = 3'b110;
        rom_memory[10985] = 3'b110;
        rom_memory[10986] = 3'b110;
        rom_memory[10987] = 3'b110;
        rom_memory[10988] = 3'b110;
        rom_memory[10989] = 3'b110;
        rom_memory[10990] = 3'b110;
        rom_memory[10991] = 3'b110;
        rom_memory[10992] = 3'b110;
        rom_memory[10993] = 3'b110;
        rom_memory[10994] = 3'b110;
        rom_memory[10995] = 3'b110;
        rom_memory[10996] = 3'b110;
        rom_memory[10997] = 3'b110;
        rom_memory[10998] = 3'b110;
        rom_memory[10999] = 3'b110;
        rom_memory[11000] = 3'b110;
        rom_memory[11001] = 3'b110;
        rom_memory[11002] = 3'b110;
        rom_memory[11003] = 3'b110;
        rom_memory[11004] = 3'b110;
        rom_memory[11005] = 3'b110;
        rom_memory[11006] = 3'b110;
        rom_memory[11007] = 3'b110;
        rom_memory[11008] = 3'b110;
        rom_memory[11009] = 3'b110;
        rom_memory[11010] = 3'b110;
        rom_memory[11011] = 3'b110;
        rom_memory[11012] = 3'b110;
        rom_memory[11013] = 3'b110;
        rom_memory[11014] = 3'b110;
        rom_memory[11015] = 3'b110;
        rom_memory[11016] = 3'b110;
        rom_memory[11017] = 3'b110;
        rom_memory[11018] = 3'b110;
        rom_memory[11019] = 3'b110;
        rom_memory[11020] = 3'b110;
        rom_memory[11021] = 3'b110;
        rom_memory[11022] = 3'b110;
        rom_memory[11023] = 3'b110;
        rom_memory[11024] = 3'b110;
        rom_memory[11025] = 3'b110;
        rom_memory[11026] = 3'b110;
        rom_memory[11027] = 3'b110;
        rom_memory[11028] = 3'b110;
        rom_memory[11029] = 3'b110;
        rom_memory[11030] = 3'b110;
        rom_memory[11031] = 3'b110;
        rom_memory[11032] = 3'b110;
        rom_memory[11033] = 3'b110;
        rom_memory[11034] = 3'b110;
        rom_memory[11035] = 3'b110;
        rom_memory[11036] = 3'b110;
        rom_memory[11037] = 3'b110;
        rom_memory[11038] = 3'b110;
        rom_memory[11039] = 3'b110;
        rom_memory[11040] = 3'b110;
        rom_memory[11041] = 3'b110;
        rom_memory[11042] = 3'b110;
        rom_memory[11043] = 3'b110;
        rom_memory[11044] = 3'b110;
        rom_memory[11045] = 3'b110;
        rom_memory[11046] = 3'b110;
        rom_memory[11047] = 3'b110;
        rom_memory[11048] = 3'b110;
        rom_memory[11049] = 3'b110;
        rom_memory[11050] = 3'b110;
        rom_memory[11051] = 3'b110;
        rom_memory[11052] = 3'b110;
        rom_memory[11053] = 3'b110;
        rom_memory[11054] = 3'b110;
        rom_memory[11055] = 3'b110;
        rom_memory[11056] = 3'b110;
        rom_memory[11057] = 3'b110;
        rom_memory[11058] = 3'b110;
        rom_memory[11059] = 3'b110;
        rom_memory[11060] = 3'b110;
        rom_memory[11061] = 3'b110;
        rom_memory[11062] = 3'b110;
        rom_memory[11063] = 3'b110;
        rom_memory[11064] = 3'b110;
        rom_memory[11065] = 3'b110;
        rom_memory[11066] = 3'b110;
        rom_memory[11067] = 3'b110;
        rom_memory[11068] = 3'b110;
        rom_memory[11069] = 3'b110;
        rom_memory[11070] = 3'b110;
        rom_memory[11071] = 3'b110;
        rom_memory[11072] = 3'b110;
        rom_memory[11073] = 3'b110;
        rom_memory[11074] = 3'b110;
        rom_memory[11075] = 3'b110;
        rom_memory[11076] = 3'b110;
        rom_memory[11077] = 3'b110;
        rom_memory[11078] = 3'b110;
        rom_memory[11079] = 3'b110;
        rom_memory[11080] = 3'b110;
        rom_memory[11081] = 3'b110;
        rom_memory[11082] = 3'b110;
        rom_memory[11083] = 3'b110;
        rom_memory[11084] = 3'b110;
        rom_memory[11085] = 3'b110;
        rom_memory[11086] = 3'b111;
        rom_memory[11087] = 3'b111;
        rom_memory[11088] = 3'b000;
        rom_memory[11089] = 3'b000;
        rom_memory[11090] = 3'b000;
        rom_memory[11091] = 3'b000;
        rom_memory[11092] = 3'b000;
        rom_memory[11093] = 3'b000;
        rom_memory[11094] = 3'b000;
        rom_memory[11095] = 3'b000;
        rom_memory[11096] = 3'b000;
        rom_memory[11097] = 3'b000;
        rom_memory[11098] = 3'b000;
        rom_memory[11099] = 3'b000;
        rom_memory[11100] = 3'b000;
        rom_memory[11101] = 3'b000;
        rom_memory[11102] = 3'b000;
        rom_memory[11103] = 3'b000;
        rom_memory[11104] = 3'b000;
        rom_memory[11105] = 3'b000;
        rom_memory[11106] = 3'b000;
        rom_memory[11107] = 3'b000;
        rom_memory[11108] = 3'b000;
        rom_memory[11109] = 3'b000;
        rom_memory[11110] = 3'b000;
        rom_memory[11111] = 3'b000;
        rom_memory[11112] = 3'b000;
        rom_memory[11113] = 3'b000;
        rom_memory[11114] = 3'b000;
        rom_memory[11115] = 3'b000;
        rom_memory[11116] = 3'b000;
        rom_memory[11117] = 3'b000;
        rom_memory[11118] = 3'b000;
        rom_memory[11119] = 3'b000;
        rom_memory[11120] = 3'b000;
        rom_memory[11121] = 3'b010;
        rom_memory[11122] = 3'b011;
        rom_memory[11123] = 3'b010;
        rom_memory[11124] = 3'b000;
        rom_memory[11125] = 3'b011;
        rom_memory[11126] = 3'b011;
        rom_memory[11127] = 3'b011;
        rom_memory[11128] = 3'b011;
        rom_memory[11129] = 3'b011;
        rom_memory[11130] = 3'b011;
        rom_memory[11131] = 3'b011;
        rom_memory[11132] = 3'b000;
        rom_memory[11133] = 3'b011;
        rom_memory[11134] = 3'b011;
        rom_memory[11135] = 3'b011;
        rom_memory[11136] = 3'b011;
        rom_memory[11137] = 3'b011;
        rom_memory[11138] = 3'b111;
        rom_memory[11139] = 3'b111;
        rom_memory[11140] = 3'b111;
        rom_memory[11141] = 3'b110;
        rom_memory[11142] = 3'b110;
        rom_memory[11143] = 3'b110;
        rom_memory[11144] = 3'b110;
        rom_memory[11145] = 3'b110;
        rom_memory[11146] = 3'b110;
        rom_memory[11147] = 3'b110;
        rom_memory[11148] = 3'b110;
        rom_memory[11149] = 3'b110;
        rom_memory[11150] = 3'b110;
        rom_memory[11151] = 3'b110;
        rom_memory[11152] = 3'b110;
        rom_memory[11153] = 3'b110;
        rom_memory[11154] = 3'b110;
        rom_memory[11155] = 3'b110;
        rom_memory[11156] = 3'b110;
        rom_memory[11157] = 3'b110;
        rom_memory[11158] = 3'b110;
        rom_memory[11159] = 3'b110;
        rom_memory[11160] = 3'b110;
        rom_memory[11161] = 3'b110;
        rom_memory[11162] = 3'b110;
        rom_memory[11163] = 3'b110;
        rom_memory[11164] = 3'b110;
        rom_memory[11165] = 3'b110;
        rom_memory[11166] = 3'b110;
        rom_memory[11167] = 3'b110;
        rom_memory[11168] = 3'b110;
        rom_memory[11169] = 3'b110;
        rom_memory[11170] = 3'b110;
        rom_memory[11171] = 3'b110;
        rom_memory[11172] = 3'b110;
        rom_memory[11173] = 3'b110;
        rom_memory[11174] = 3'b110;
        rom_memory[11175] = 3'b110;
        rom_memory[11176] = 3'b110;
        rom_memory[11177] = 3'b110;
        rom_memory[11178] = 3'b110;
        rom_memory[11179] = 3'b110;
        rom_memory[11180] = 3'b110;
        rom_memory[11181] = 3'b110;
        rom_memory[11182] = 3'b110;
        rom_memory[11183] = 3'b110;
        rom_memory[11184] = 3'b110;
        rom_memory[11185] = 3'b110;
        rom_memory[11186] = 3'b110;
        rom_memory[11187] = 3'b110;
        rom_memory[11188] = 3'b110;
        rom_memory[11189] = 3'b110;
        rom_memory[11190] = 3'b110;
        rom_memory[11191] = 3'b110;
        rom_memory[11192] = 3'b110;
        rom_memory[11193] = 3'b110;
        rom_memory[11194] = 3'b110;
        rom_memory[11195] = 3'b110;
        rom_memory[11196] = 3'b110;
        rom_memory[11197] = 3'b110;
        rom_memory[11198] = 3'b110;
        rom_memory[11199] = 3'b110;
        rom_memory[11200] = 3'b110;
        rom_memory[11201] = 3'b110;
        rom_memory[11202] = 3'b110;
        rom_memory[11203] = 3'b110;
        rom_memory[11204] = 3'b110;
        rom_memory[11205] = 3'b110;
        rom_memory[11206] = 3'b110;
        rom_memory[11207] = 3'b110;
        rom_memory[11208] = 3'b110;
        rom_memory[11209] = 3'b110;
        rom_memory[11210] = 3'b110;
        rom_memory[11211] = 3'b110;
        rom_memory[11212] = 3'b110;
        rom_memory[11213] = 3'b110;
        rom_memory[11214] = 3'b110;
        rom_memory[11215] = 3'b110;
        rom_memory[11216] = 3'b110;
        rom_memory[11217] = 3'b110;
        rom_memory[11218] = 3'b110;
        rom_memory[11219] = 3'b110;
        rom_memory[11220] = 3'b110;
        rom_memory[11221] = 3'b110;
        rom_memory[11222] = 3'b110;
        rom_memory[11223] = 3'b110;
        rom_memory[11224] = 3'b110;
        rom_memory[11225] = 3'b110;
        rom_memory[11226] = 3'b110;
        rom_memory[11227] = 3'b110;
        rom_memory[11228] = 3'b110;
        rom_memory[11229] = 3'b110;
        rom_memory[11230] = 3'b110;
        rom_memory[11231] = 3'b110;
        rom_memory[11232] = 3'b110;
        rom_memory[11233] = 3'b110;
        rom_memory[11234] = 3'b110;
        rom_memory[11235] = 3'b110;
        rom_memory[11236] = 3'b110;
        rom_memory[11237] = 3'b110;
        rom_memory[11238] = 3'b110;
        rom_memory[11239] = 3'b110;
        rom_memory[11240] = 3'b110;
        rom_memory[11241] = 3'b110;
        rom_memory[11242] = 3'b110;
        rom_memory[11243] = 3'b110;
        rom_memory[11244] = 3'b110;
        rom_memory[11245] = 3'b110;
        rom_memory[11246] = 3'b110;
        rom_memory[11247] = 3'b110;
        rom_memory[11248] = 3'b110;
        rom_memory[11249] = 3'b110;
        rom_memory[11250] = 3'b110;
        rom_memory[11251] = 3'b110;
        rom_memory[11252] = 3'b110;
        rom_memory[11253] = 3'b110;
        rom_memory[11254] = 3'b110;
        rom_memory[11255] = 3'b110;
        rom_memory[11256] = 3'b110;
        rom_memory[11257] = 3'b110;
        rom_memory[11258] = 3'b110;
        rom_memory[11259] = 3'b110;
        rom_memory[11260] = 3'b110;
        rom_memory[11261] = 3'b110;
        rom_memory[11262] = 3'b110;
        rom_memory[11263] = 3'b110;
        rom_memory[11264] = 3'b110;
        rom_memory[11265] = 3'b110;
        rom_memory[11266] = 3'b110;
        rom_memory[11267] = 3'b110;
        rom_memory[11268] = 3'b110;
        rom_memory[11269] = 3'b110;
        rom_memory[11270] = 3'b110;
        rom_memory[11271] = 3'b110;
        rom_memory[11272] = 3'b110;
        rom_memory[11273] = 3'b110;
        rom_memory[11274] = 3'b110;
        rom_memory[11275] = 3'b110;
        rom_memory[11276] = 3'b110;
        rom_memory[11277] = 3'b110;
        rom_memory[11278] = 3'b110;
        rom_memory[11279] = 3'b110;
        rom_memory[11280] = 3'b110;
        rom_memory[11281] = 3'b110;
        rom_memory[11282] = 3'b110;
        rom_memory[11283] = 3'b110;
        rom_memory[11284] = 3'b110;
        rom_memory[11285] = 3'b110;
        rom_memory[11286] = 3'b110;
        rom_memory[11287] = 3'b110;
        rom_memory[11288] = 3'b110;
        rom_memory[11289] = 3'b110;
        rom_memory[11290] = 3'b110;
        rom_memory[11291] = 3'b110;
        rom_memory[11292] = 3'b110;
        rom_memory[11293] = 3'b110;
        rom_memory[11294] = 3'b110;
        rom_memory[11295] = 3'b110;
        rom_memory[11296] = 3'b110;
        rom_memory[11297] = 3'b110;
        rom_memory[11298] = 3'b110;
        rom_memory[11299] = 3'b110;
        rom_memory[11300] = 3'b110;
        rom_memory[11301] = 3'b110;
        rom_memory[11302] = 3'b110;
        rom_memory[11303] = 3'b110;
        rom_memory[11304] = 3'b110;
        rom_memory[11305] = 3'b110;
        rom_memory[11306] = 3'b110;
        rom_memory[11307] = 3'b110;
        rom_memory[11308] = 3'b110;
        rom_memory[11309] = 3'b110;
        rom_memory[11310] = 3'b110;
        rom_memory[11311] = 3'b110;
        rom_memory[11312] = 3'b110;
        rom_memory[11313] = 3'b110;
        rom_memory[11314] = 3'b110;
        rom_memory[11315] = 3'b110;
        rom_memory[11316] = 3'b110;
        rom_memory[11317] = 3'b110;
        rom_memory[11318] = 3'b110;
        rom_memory[11319] = 3'b110;
        rom_memory[11320] = 3'b110;
        rom_memory[11321] = 3'b110;
        rom_memory[11322] = 3'b110;
        rom_memory[11323] = 3'b110;
        rom_memory[11324] = 3'b110;
        rom_memory[11325] = 3'b110;
        rom_memory[11326] = 3'b110;
        rom_memory[11327] = 3'b111;
        rom_memory[11328] = 3'b000;
        rom_memory[11329] = 3'b000;
        rom_memory[11330] = 3'b000;
        rom_memory[11331] = 3'b000;
        rom_memory[11332] = 3'b000;
        rom_memory[11333] = 3'b000;
        rom_memory[11334] = 3'b000;
        rom_memory[11335] = 3'b000;
        rom_memory[11336] = 3'b000;
        rom_memory[11337] = 3'b000;
        rom_memory[11338] = 3'b000;
        rom_memory[11339] = 3'b000;
        rom_memory[11340] = 3'b000;
        rom_memory[11341] = 3'b000;
        rom_memory[11342] = 3'b000;
        rom_memory[11343] = 3'b000;
        rom_memory[11344] = 3'b000;
        rom_memory[11345] = 3'b000;
        rom_memory[11346] = 3'b000;
        rom_memory[11347] = 3'b000;
        rom_memory[11348] = 3'b000;
        rom_memory[11349] = 3'b000;
        rom_memory[11350] = 3'b000;
        rom_memory[11351] = 3'b000;
        rom_memory[11352] = 3'b000;
        rom_memory[11353] = 3'b000;
        rom_memory[11354] = 3'b000;
        rom_memory[11355] = 3'b000;
        rom_memory[11356] = 3'b000;
        rom_memory[11357] = 3'b000;
        rom_memory[11358] = 3'b000;
        rom_memory[11359] = 3'b000;
        rom_memory[11360] = 3'b000;
        rom_memory[11361] = 3'b011;
        rom_memory[11362] = 3'b011;
        rom_memory[11363] = 3'b000;
        rom_memory[11364] = 3'b010;
        rom_memory[11365] = 3'b011;
        rom_memory[11366] = 3'b010;
        rom_memory[11367] = 3'b011;
        rom_memory[11368] = 3'b011;
        rom_memory[11369] = 3'b011;
        rom_memory[11370] = 3'b011;
        rom_memory[11371] = 3'b011;
        rom_memory[11372] = 3'b001;
        rom_memory[11373] = 3'b011;
        rom_memory[11374] = 3'b011;
        rom_memory[11375] = 3'b011;
        rom_memory[11376] = 3'b011;
        rom_memory[11377] = 3'b001;
        rom_memory[11378] = 3'b011;
        rom_memory[11379] = 3'b111;
        rom_memory[11380] = 3'b111;
        rom_memory[11381] = 3'b111;
        rom_memory[11382] = 3'b110;
        rom_memory[11383] = 3'b110;
        rom_memory[11384] = 3'b110;
        rom_memory[11385] = 3'b110;
        rom_memory[11386] = 3'b110;
        rom_memory[11387] = 3'b110;
        rom_memory[11388] = 3'b110;
        rom_memory[11389] = 3'b110;
        rom_memory[11390] = 3'b110;
        rom_memory[11391] = 3'b110;
        rom_memory[11392] = 3'b110;
        rom_memory[11393] = 3'b110;
        rom_memory[11394] = 3'b110;
        rom_memory[11395] = 3'b110;
        rom_memory[11396] = 3'b110;
        rom_memory[11397] = 3'b110;
        rom_memory[11398] = 3'b110;
        rom_memory[11399] = 3'b110;
        rom_memory[11400] = 3'b110;
        rom_memory[11401] = 3'b110;
        rom_memory[11402] = 3'b110;
        rom_memory[11403] = 3'b110;
        rom_memory[11404] = 3'b110;
        rom_memory[11405] = 3'b110;
        rom_memory[11406] = 3'b110;
        rom_memory[11407] = 3'b110;
        rom_memory[11408] = 3'b110;
        rom_memory[11409] = 3'b110;
        rom_memory[11410] = 3'b110;
        rom_memory[11411] = 3'b110;
        rom_memory[11412] = 3'b110;
        rom_memory[11413] = 3'b110;
        rom_memory[11414] = 3'b110;
        rom_memory[11415] = 3'b110;
        rom_memory[11416] = 3'b110;
        rom_memory[11417] = 3'b110;
        rom_memory[11418] = 3'b110;
        rom_memory[11419] = 3'b110;
        rom_memory[11420] = 3'b110;
        rom_memory[11421] = 3'b110;
        rom_memory[11422] = 3'b110;
        rom_memory[11423] = 3'b110;
        rom_memory[11424] = 3'b110;
        rom_memory[11425] = 3'b110;
        rom_memory[11426] = 3'b110;
        rom_memory[11427] = 3'b110;
        rom_memory[11428] = 3'b110;
        rom_memory[11429] = 3'b110;
        rom_memory[11430] = 3'b110;
        rom_memory[11431] = 3'b110;
        rom_memory[11432] = 3'b110;
        rom_memory[11433] = 3'b110;
        rom_memory[11434] = 3'b110;
        rom_memory[11435] = 3'b110;
        rom_memory[11436] = 3'b110;
        rom_memory[11437] = 3'b110;
        rom_memory[11438] = 3'b110;
        rom_memory[11439] = 3'b110;
        rom_memory[11440] = 3'b110;
        rom_memory[11441] = 3'b110;
        rom_memory[11442] = 3'b110;
        rom_memory[11443] = 3'b110;
        rom_memory[11444] = 3'b110;
        rom_memory[11445] = 3'b110;
        rom_memory[11446] = 3'b110;
        rom_memory[11447] = 3'b110;
        rom_memory[11448] = 3'b110;
        rom_memory[11449] = 3'b110;
        rom_memory[11450] = 3'b110;
        rom_memory[11451] = 3'b110;
        rom_memory[11452] = 3'b110;
        rom_memory[11453] = 3'b110;
        rom_memory[11454] = 3'b110;
        rom_memory[11455] = 3'b110;
        rom_memory[11456] = 3'b110;
        rom_memory[11457] = 3'b110;
        rom_memory[11458] = 3'b110;
        rom_memory[11459] = 3'b110;
        rom_memory[11460] = 3'b110;
        rom_memory[11461] = 3'b110;
        rom_memory[11462] = 3'b110;
        rom_memory[11463] = 3'b110;
        rom_memory[11464] = 3'b110;
        rom_memory[11465] = 3'b110;
        rom_memory[11466] = 3'b110;
        rom_memory[11467] = 3'b110;
        rom_memory[11468] = 3'b110;
        rom_memory[11469] = 3'b110;
        rom_memory[11470] = 3'b110;
        rom_memory[11471] = 3'b110;
        rom_memory[11472] = 3'b110;
        rom_memory[11473] = 3'b110;
        rom_memory[11474] = 3'b110;
        rom_memory[11475] = 3'b110;
        rom_memory[11476] = 3'b110;
        rom_memory[11477] = 3'b110;
        rom_memory[11478] = 3'b110;
        rom_memory[11479] = 3'b110;
        rom_memory[11480] = 3'b110;
        rom_memory[11481] = 3'b110;
        rom_memory[11482] = 3'b110;
        rom_memory[11483] = 3'b110;
        rom_memory[11484] = 3'b110;
        rom_memory[11485] = 3'b110;
        rom_memory[11486] = 3'b110;
        rom_memory[11487] = 3'b110;
        rom_memory[11488] = 3'b110;
        rom_memory[11489] = 3'b110;
        rom_memory[11490] = 3'b110;
        rom_memory[11491] = 3'b110;
        rom_memory[11492] = 3'b110;
        rom_memory[11493] = 3'b110;
        rom_memory[11494] = 3'b110;
        rom_memory[11495] = 3'b110;
        rom_memory[11496] = 3'b110;
        rom_memory[11497] = 3'b110;
        rom_memory[11498] = 3'b110;
        rom_memory[11499] = 3'b110;
        rom_memory[11500] = 3'b110;
        rom_memory[11501] = 3'b110;
        rom_memory[11502] = 3'b110;
        rom_memory[11503] = 3'b110;
        rom_memory[11504] = 3'b110;
        rom_memory[11505] = 3'b110;
        rom_memory[11506] = 3'b110;
        rom_memory[11507] = 3'b110;
        rom_memory[11508] = 3'b110;
        rom_memory[11509] = 3'b110;
        rom_memory[11510] = 3'b110;
        rom_memory[11511] = 3'b110;
        rom_memory[11512] = 3'b110;
        rom_memory[11513] = 3'b110;
        rom_memory[11514] = 3'b110;
        rom_memory[11515] = 3'b110;
        rom_memory[11516] = 3'b110;
        rom_memory[11517] = 3'b110;
        rom_memory[11518] = 3'b110;
        rom_memory[11519] = 3'b110;
        rom_memory[11520] = 3'b110;
        rom_memory[11521] = 3'b110;
        rom_memory[11522] = 3'b110;
        rom_memory[11523] = 3'b110;
        rom_memory[11524] = 3'b110;
        rom_memory[11525] = 3'b110;
        rom_memory[11526] = 3'b110;
        rom_memory[11527] = 3'b110;
        rom_memory[11528] = 3'b110;
        rom_memory[11529] = 3'b110;
        rom_memory[11530] = 3'b110;
        rom_memory[11531] = 3'b110;
        rom_memory[11532] = 3'b110;
        rom_memory[11533] = 3'b110;
        rom_memory[11534] = 3'b110;
        rom_memory[11535] = 3'b110;
        rom_memory[11536] = 3'b110;
        rom_memory[11537] = 3'b110;
        rom_memory[11538] = 3'b110;
        rom_memory[11539] = 3'b110;
        rom_memory[11540] = 3'b110;
        rom_memory[11541] = 3'b110;
        rom_memory[11542] = 3'b110;
        rom_memory[11543] = 3'b110;
        rom_memory[11544] = 3'b110;
        rom_memory[11545] = 3'b110;
        rom_memory[11546] = 3'b110;
        rom_memory[11547] = 3'b110;
        rom_memory[11548] = 3'b110;
        rom_memory[11549] = 3'b110;
        rom_memory[11550] = 3'b110;
        rom_memory[11551] = 3'b110;
        rom_memory[11552] = 3'b110;
        rom_memory[11553] = 3'b110;
        rom_memory[11554] = 3'b110;
        rom_memory[11555] = 3'b110;
        rom_memory[11556] = 3'b110;
        rom_memory[11557] = 3'b110;
        rom_memory[11558] = 3'b110;
        rom_memory[11559] = 3'b110;
        rom_memory[11560] = 3'b110;
        rom_memory[11561] = 3'b110;
        rom_memory[11562] = 3'b110;
        rom_memory[11563] = 3'b110;
        rom_memory[11564] = 3'b110;
        rom_memory[11565] = 3'b110;
        rom_memory[11566] = 3'b110;
        rom_memory[11567] = 3'b111;
        rom_memory[11568] = 3'b000;
        rom_memory[11569] = 3'b000;
        rom_memory[11570] = 3'b000;
        rom_memory[11571] = 3'b000;
        rom_memory[11572] = 3'b000;
        rom_memory[11573] = 3'b000;
        rom_memory[11574] = 3'b000;
        rom_memory[11575] = 3'b000;
        rom_memory[11576] = 3'b000;
        rom_memory[11577] = 3'b000;
        rom_memory[11578] = 3'b000;
        rom_memory[11579] = 3'b000;
        rom_memory[11580] = 3'b000;
        rom_memory[11581] = 3'b000;
        rom_memory[11582] = 3'b000;
        rom_memory[11583] = 3'b000;
        rom_memory[11584] = 3'b000;
        rom_memory[11585] = 3'b000;
        rom_memory[11586] = 3'b000;
        rom_memory[11587] = 3'b000;
        rom_memory[11588] = 3'b000;
        rom_memory[11589] = 3'b000;
        rom_memory[11590] = 3'b000;
        rom_memory[11591] = 3'b000;
        rom_memory[11592] = 3'b000;
        rom_memory[11593] = 3'b000;
        rom_memory[11594] = 3'b000;
        rom_memory[11595] = 3'b000;
        rom_memory[11596] = 3'b000;
        rom_memory[11597] = 3'b000;
        rom_memory[11598] = 3'b000;
        rom_memory[11599] = 3'b000;
        rom_memory[11600] = 3'b000;
        rom_memory[11601] = 3'b000;
        rom_memory[11602] = 3'b000;
        rom_memory[11603] = 3'b000;
        rom_memory[11604] = 3'b000;
        rom_memory[11605] = 3'b000;
        rom_memory[11606] = 3'b000;
        rom_memory[11607] = 3'b000;
        rom_memory[11608] = 3'b000;
        rom_memory[11609] = 3'b010;
        rom_memory[11610] = 3'b011;
        rom_memory[11611] = 3'b011;
        rom_memory[11612] = 3'b011;
        rom_memory[11613] = 3'b000;
        rom_memory[11614] = 3'b011;
        rom_memory[11615] = 3'b011;
        rom_memory[11616] = 3'b011;
        rom_memory[11617] = 3'b011;
        rom_memory[11618] = 3'b011;
        rom_memory[11619] = 3'b011;
        rom_memory[11620] = 3'b001;
        rom_memory[11621] = 3'b111;
        rom_memory[11622] = 3'b110;
        rom_memory[11623] = 3'b110;
        rom_memory[11624] = 3'b111;
        rom_memory[11625] = 3'b110;
        rom_memory[11626] = 3'b110;
        rom_memory[11627] = 3'b110;
        rom_memory[11628] = 3'b110;
        rom_memory[11629] = 3'b110;
        rom_memory[11630] = 3'b110;
        rom_memory[11631] = 3'b110;
        rom_memory[11632] = 3'b110;
        rom_memory[11633] = 3'b110;
        rom_memory[11634] = 3'b110;
        rom_memory[11635] = 3'b110;
        rom_memory[11636] = 3'b110;
        rom_memory[11637] = 3'b110;
        rom_memory[11638] = 3'b110;
        rom_memory[11639] = 3'b110;
        rom_memory[11640] = 3'b110;
        rom_memory[11641] = 3'b110;
        rom_memory[11642] = 3'b110;
        rom_memory[11643] = 3'b110;
        rom_memory[11644] = 3'b110;
        rom_memory[11645] = 3'b110;
        rom_memory[11646] = 3'b110;
        rom_memory[11647] = 3'b110;
        rom_memory[11648] = 3'b110;
        rom_memory[11649] = 3'b110;
        rom_memory[11650] = 3'b110;
        rom_memory[11651] = 3'b110;
        rom_memory[11652] = 3'b110;
        rom_memory[11653] = 3'b110;
        rom_memory[11654] = 3'b110;
        rom_memory[11655] = 3'b110;
        rom_memory[11656] = 3'b110;
        rom_memory[11657] = 3'b110;
        rom_memory[11658] = 3'b110;
        rom_memory[11659] = 3'b110;
        rom_memory[11660] = 3'b110;
        rom_memory[11661] = 3'b110;
        rom_memory[11662] = 3'b110;
        rom_memory[11663] = 3'b110;
        rom_memory[11664] = 3'b110;
        rom_memory[11665] = 3'b110;
        rom_memory[11666] = 3'b110;
        rom_memory[11667] = 3'b110;
        rom_memory[11668] = 3'b110;
        rom_memory[11669] = 3'b110;
        rom_memory[11670] = 3'b110;
        rom_memory[11671] = 3'b110;
        rom_memory[11672] = 3'b110;
        rom_memory[11673] = 3'b110;
        rom_memory[11674] = 3'b110;
        rom_memory[11675] = 3'b110;
        rom_memory[11676] = 3'b110;
        rom_memory[11677] = 3'b110;
        rom_memory[11678] = 3'b110;
        rom_memory[11679] = 3'b110;
        rom_memory[11680] = 3'b110;
        rom_memory[11681] = 3'b110;
        rom_memory[11682] = 3'b110;
        rom_memory[11683] = 3'b110;
        rom_memory[11684] = 3'b110;
        rom_memory[11685] = 3'b110;
        rom_memory[11686] = 3'b110;
        rom_memory[11687] = 3'b110;
        rom_memory[11688] = 3'b110;
        rom_memory[11689] = 3'b110;
        rom_memory[11690] = 3'b110;
        rom_memory[11691] = 3'b110;
        rom_memory[11692] = 3'b110;
        rom_memory[11693] = 3'b110;
        rom_memory[11694] = 3'b110;
        rom_memory[11695] = 3'b110;
        rom_memory[11696] = 3'b110;
        rom_memory[11697] = 3'b110;
        rom_memory[11698] = 3'b110;
        rom_memory[11699] = 3'b110;
        rom_memory[11700] = 3'b110;
        rom_memory[11701] = 3'b110;
        rom_memory[11702] = 3'b110;
        rom_memory[11703] = 3'b110;
        rom_memory[11704] = 3'b110;
        rom_memory[11705] = 3'b110;
        rom_memory[11706] = 3'b110;
        rom_memory[11707] = 3'b110;
        rom_memory[11708] = 3'b110;
        rom_memory[11709] = 3'b110;
        rom_memory[11710] = 3'b110;
        rom_memory[11711] = 3'b110;
        rom_memory[11712] = 3'b110;
        rom_memory[11713] = 3'b110;
        rom_memory[11714] = 3'b110;
        rom_memory[11715] = 3'b110;
        rom_memory[11716] = 3'b110;
        rom_memory[11717] = 3'b110;
        rom_memory[11718] = 3'b110;
        rom_memory[11719] = 3'b110;
        rom_memory[11720] = 3'b110;
        rom_memory[11721] = 3'b110;
        rom_memory[11722] = 3'b110;
        rom_memory[11723] = 3'b110;
        rom_memory[11724] = 3'b110;
        rom_memory[11725] = 3'b110;
        rom_memory[11726] = 3'b110;
        rom_memory[11727] = 3'b110;
        rom_memory[11728] = 3'b110;
        rom_memory[11729] = 3'b110;
        rom_memory[11730] = 3'b110;
        rom_memory[11731] = 3'b110;
        rom_memory[11732] = 3'b110;
        rom_memory[11733] = 3'b110;
        rom_memory[11734] = 3'b110;
        rom_memory[11735] = 3'b110;
        rom_memory[11736] = 3'b110;
        rom_memory[11737] = 3'b110;
        rom_memory[11738] = 3'b110;
        rom_memory[11739] = 3'b110;
        rom_memory[11740] = 3'b110;
        rom_memory[11741] = 3'b110;
        rom_memory[11742] = 3'b110;
        rom_memory[11743] = 3'b110;
        rom_memory[11744] = 3'b110;
        rom_memory[11745] = 3'b110;
        rom_memory[11746] = 3'b110;
        rom_memory[11747] = 3'b110;
        rom_memory[11748] = 3'b110;
        rom_memory[11749] = 3'b110;
        rom_memory[11750] = 3'b110;
        rom_memory[11751] = 3'b110;
        rom_memory[11752] = 3'b110;
        rom_memory[11753] = 3'b110;
        rom_memory[11754] = 3'b110;
        rom_memory[11755] = 3'b110;
        rom_memory[11756] = 3'b110;
        rom_memory[11757] = 3'b110;
        rom_memory[11758] = 3'b110;
        rom_memory[11759] = 3'b110;
        rom_memory[11760] = 3'b110;
        rom_memory[11761] = 3'b110;
        rom_memory[11762] = 3'b110;
        rom_memory[11763] = 3'b110;
        rom_memory[11764] = 3'b110;
        rom_memory[11765] = 3'b110;
        rom_memory[11766] = 3'b110;
        rom_memory[11767] = 3'b110;
        rom_memory[11768] = 3'b110;
        rom_memory[11769] = 3'b110;
        rom_memory[11770] = 3'b110;
        rom_memory[11771] = 3'b110;
        rom_memory[11772] = 3'b110;
        rom_memory[11773] = 3'b110;
        rom_memory[11774] = 3'b110;
        rom_memory[11775] = 3'b110;
        rom_memory[11776] = 3'b110;
        rom_memory[11777] = 3'b110;
        rom_memory[11778] = 3'b110;
        rom_memory[11779] = 3'b110;
        rom_memory[11780] = 3'b110;
        rom_memory[11781] = 3'b110;
        rom_memory[11782] = 3'b110;
        rom_memory[11783] = 3'b110;
        rom_memory[11784] = 3'b110;
        rom_memory[11785] = 3'b110;
        rom_memory[11786] = 3'b110;
        rom_memory[11787] = 3'b110;
        rom_memory[11788] = 3'b110;
        rom_memory[11789] = 3'b110;
        rom_memory[11790] = 3'b110;
        rom_memory[11791] = 3'b110;
        rom_memory[11792] = 3'b110;
        rom_memory[11793] = 3'b110;
        rom_memory[11794] = 3'b110;
        rom_memory[11795] = 3'b110;
        rom_memory[11796] = 3'b110;
        rom_memory[11797] = 3'b110;
        rom_memory[11798] = 3'b110;
        rom_memory[11799] = 3'b110;
        rom_memory[11800] = 3'b110;
        rom_memory[11801] = 3'b110;
        rom_memory[11802] = 3'b110;
        rom_memory[11803] = 3'b110;
        rom_memory[11804] = 3'b110;
        rom_memory[11805] = 3'b110;
        rom_memory[11806] = 3'b111;
        rom_memory[11807] = 3'b111;
        rom_memory[11808] = 3'b000;
        rom_memory[11809] = 3'b000;
        rom_memory[11810] = 3'b000;
        rom_memory[11811] = 3'b000;
        rom_memory[11812] = 3'b000;
        rom_memory[11813] = 3'b000;
        rom_memory[11814] = 3'b000;
        rom_memory[11815] = 3'b000;
        rom_memory[11816] = 3'b000;
        rom_memory[11817] = 3'b000;
        rom_memory[11818] = 3'b000;
        rom_memory[11819] = 3'b000;
        rom_memory[11820] = 3'b000;
        rom_memory[11821] = 3'b000;
        rom_memory[11822] = 3'b000;
        rom_memory[11823] = 3'b000;
        rom_memory[11824] = 3'b000;
        rom_memory[11825] = 3'b000;
        rom_memory[11826] = 3'b000;
        rom_memory[11827] = 3'b000;
        rom_memory[11828] = 3'b000;
        rom_memory[11829] = 3'b000;
        rom_memory[11830] = 3'b000;
        rom_memory[11831] = 3'b000;
        rom_memory[11832] = 3'b000;
        rom_memory[11833] = 3'b000;
        rom_memory[11834] = 3'b000;
        rom_memory[11835] = 3'b000;
        rom_memory[11836] = 3'b000;
        rom_memory[11837] = 3'b000;
        rom_memory[11838] = 3'b000;
        rom_memory[11839] = 3'b000;
        rom_memory[11840] = 3'b000;
        rom_memory[11841] = 3'b000;
        rom_memory[11842] = 3'b000;
        rom_memory[11843] = 3'b000;
        rom_memory[11844] = 3'b000;
        rom_memory[11845] = 3'b000;
        rom_memory[11846] = 3'b011;
        rom_memory[11847] = 3'b000;
        rom_memory[11848] = 3'b010;
        rom_memory[11849] = 3'b011;
        rom_memory[11850] = 3'b011;
        rom_memory[11851] = 3'b011;
        rom_memory[11852] = 3'b000;
        rom_memory[11853] = 3'b000;
        rom_memory[11854] = 3'b011;
        rom_memory[11855] = 3'b011;
        rom_memory[11856] = 3'b011;
        rom_memory[11857] = 3'b011;
        rom_memory[11858] = 3'b011;
        rom_memory[11859] = 3'b011;
        rom_memory[11860] = 3'b000;
        rom_memory[11861] = 3'b111;
        rom_memory[11862] = 3'b111;
        rom_memory[11863] = 3'b111;
        rom_memory[11864] = 3'b111;
        rom_memory[11865] = 3'b110;
        rom_memory[11866] = 3'b110;
        rom_memory[11867] = 3'b110;
        rom_memory[11868] = 3'b110;
        rom_memory[11869] = 3'b110;
        rom_memory[11870] = 3'b110;
        rom_memory[11871] = 3'b110;
        rom_memory[11872] = 3'b110;
        rom_memory[11873] = 3'b110;
        rom_memory[11874] = 3'b110;
        rom_memory[11875] = 3'b110;
        rom_memory[11876] = 3'b110;
        rom_memory[11877] = 3'b110;
        rom_memory[11878] = 3'b110;
        rom_memory[11879] = 3'b110;
        rom_memory[11880] = 3'b110;
        rom_memory[11881] = 3'b110;
        rom_memory[11882] = 3'b110;
        rom_memory[11883] = 3'b110;
        rom_memory[11884] = 3'b110;
        rom_memory[11885] = 3'b110;
        rom_memory[11886] = 3'b110;
        rom_memory[11887] = 3'b110;
        rom_memory[11888] = 3'b110;
        rom_memory[11889] = 3'b110;
        rom_memory[11890] = 3'b110;
        rom_memory[11891] = 3'b110;
        rom_memory[11892] = 3'b110;
        rom_memory[11893] = 3'b110;
        rom_memory[11894] = 3'b110;
        rom_memory[11895] = 3'b110;
        rom_memory[11896] = 3'b110;
        rom_memory[11897] = 3'b110;
        rom_memory[11898] = 3'b110;
        rom_memory[11899] = 3'b110;
        rom_memory[11900] = 3'b110;
        rom_memory[11901] = 3'b110;
        rom_memory[11902] = 3'b110;
        rom_memory[11903] = 3'b110;
        rom_memory[11904] = 3'b110;
        rom_memory[11905] = 3'b110;
        rom_memory[11906] = 3'b110;
        rom_memory[11907] = 3'b110;
        rom_memory[11908] = 3'b110;
        rom_memory[11909] = 3'b110;
        rom_memory[11910] = 3'b110;
        rom_memory[11911] = 3'b110;
        rom_memory[11912] = 3'b110;
        rom_memory[11913] = 3'b110;
        rom_memory[11914] = 3'b110;
        rom_memory[11915] = 3'b110;
        rom_memory[11916] = 3'b110;
        rom_memory[11917] = 3'b110;
        rom_memory[11918] = 3'b110;
        rom_memory[11919] = 3'b110;
        rom_memory[11920] = 3'b110;
        rom_memory[11921] = 3'b110;
        rom_memory[11922] = 3'b110;
        rom_memory[11923] = 3'b110;
        rom_memory[11924] = 3'b110;
        rom_memory[11925] = 3'b110;
        rom_memory[11926] = 3'b110;
        rom_memory[11927] = 3'b110;
        rom_memory[11928] = 3'b110;
        rom_memory[11929] = 3'b110;
        rom_memory[11930] = 3'b110;
        rom_memory[11931] = 3'b110;
        rom_memory[11932] = 3'b110;
        rom_memory[11933] = 3'b110;
        rom_memory[11934] = 3'b110;
        rom_memory[11935] = 3'b110;
        rom_memory[11936] = 3'b110;
        rom_memory[11937] = 3'b110;
        rom_memory[11938] = 3'b110;
        rom_memory[11939] = 3'b110;
        rom_memory[11940] = 3'b110;
        rom_memory[11941] = 3'b110;
        rom_memory[11942] = 3'b110;
        rom_memory[11943] = 3'b110;
        rom_memory[11944] = 3'b110;
        rom_memory[11945] = 3'b110;
        rom_memory[11946] = 3'b110;
        rom_memory[11947] = 3'b110;
        rom_memory[11948] = 3'b110;
        rom_memory[11949] = 3'b110;
        rom_memory[11950] = 3'b110;
        rom_memory[11951] = 3'b110;
        rom_memory[11952] = 3'b110;
        rom_memory[11953] = 3'b110;
        rom_memory[11954] = 3'b110;
        rom_memory[11955] = 3'b110;
        rom_memory[11956] = 3'b110;
        rom_memory[11957] = 3'b110;
        rom_memory[11958] = 3'b110;
        rom_memory[11959] = 3'b110;
        rom_memory[11960] = 3'b110;
        rom_memory[11961] = 3'b110;
        rom_memory[11962] = 3'b110;
        rom_memory[11963] = 3'b110;
        rom_memory[11964] = 3'b110;
        rom_memory[11965] = 3'b110;
        rom_memory[11966] = 3'b110;
        rom_memory[11967] = 3'b110;
        rom_memory[11968] = 3'b110;
        rom_memory[11969] = 3'b110;
        rom_memory[11970] = 3'b110;
        rom_memory[11971] = 3'b110;
        rom_memory[11972] = 3'b110;
        rom_memory[11973] = 3'b110;
        rom_memory[11974] = 3'b110;
        rom_memory[11975] = 3'b110;
        rom_memory[11976] = 3'b110;
        rom_memory[11977] = 3'b110;
        rom_memory[11978] = 3'b110;
        rom_memory[11979] = 3'b110;
        rom_memory[11980] = 3'b110;
        rom_memory[11981] = 3'b110;
        rom_memory[11982] = 3'b110;
        rom_memory[11983] = 3'b110;
        rom_memory[11984] = 3'b110;
        rom_memory[11985] = 3'b110;
        rom_memory[11986] = 3'b110;
        rom_memory[11987] = 3'b110;
        rom_memory[11988] = 3'b110;
        rom_memory[11989] = 3'b110;
        rom_memory[11990] = 3'b110;
        rom_memory[11991] = 3'b110;
        rom_memory[11992] = 3'b110;
        rom_memory[11993] = 3'b110;
        rom_memory[11994] = 3'b110;
        rom_memory[11995] = 3'b110;
        rom_memory[11996] = 3'b110;
        rom_memory[11997] = 3'b110;
        rom_memory[11998] = 3'b110;
        rom_memory[11999] = 3'b110;
        rom_memory[12000] = 3'b110;
        rom_memory[12001] = 3'b110;
        rom_memory[12002] = 3'b110;
        rom_memory[12003] = 3'b110;
        rom_memory[12004] = 3'b110;
        rom_memory[12005] = 3'b110;
        rom_memory[12006] = 3'b110;
        rom_memory[12007] = 3'b110;
        rom_memory[12008] = 3'b110;
        rom_memory[12009] = 3'b110;
        rom_memory[12010] = 3'b110;
        rom_memory[12011] = 3'b110;
        rom_memory[12012] = 3'b110;
        rom_memory[12013] = 3'b110;
        rom_memory[12014] = 3'b110;
        rom_memory[12015] = 3'b110;
        rom_memory[12016] = 3'b110;
        rom_memory[12017] = 3'b110;
        rom_memory[12018] = 3'b110;
        rom_memory[12019] = 3'b110;
        rom_memory[12020] = 3'b110;
        rom_memory[12021] = 3'b110;
        rom_memory[12022] = 3'b110;
        rom_memory[12023] = 3'b110;
        rom_memory[12024] = 3'b110;
        rom_memory[12025] = 3'b110;
        rom_memory[12026] = 3'b110;
        rom_memory[12027] = 3'b110;
        rom_memory[12028] = 3'b110;
        rom_memory[12029] = 3'b110;
        rom_memory[12030] = 3'b110;
        rom_memory[12031] = 3'b110;
        rom_memory[12032] = 3'b110;
        rom_memory[12033] = 3'b110;
        rom_memory[12034] = 3'b110;
        rom_memory[12035] = 3'b110;
        rom_memory[12036] = 3'b110;
        rom_memory[12037] = 3'b110;
        rom_memory[12038] = 3'b110;
        rom_memory[12039] = 3'b110;
        rom_memory[12040] = 3'b110;
        rom_memory[12041] = 3'b110;
        rom_memory[12042] = 3'b110;
        rom_memory[12043] = 3'b110;
        rom_memory[12044] = 3'b110;
        rom_memory[12045] = 3'b110;
        rom_memory[12046] = 3'b111;
        rom_memory[12047] = 3'b111;
        rom_memory[12048] = 3'b000;
        rom_memory[12049] = 3'b000;
        rom_memory[12050] = 3'b000;
        rom_memory[12051] = 3'b000;
        rom_memory[12052] = 3'b000;
        rom_memory[12053] = 3'b000;
        rom_memory[12054] = 3'b000;
        rom_memory[12055] = 3'b000;
        rom_memory[12056] = 3'b000;
        rom_memory[12057] = 3'b000;
        rom_memory[12058] = 3'b000;
        rom_memory[12059] = 3'b000;
        rom_memory[12060] = 3'b000;
        rom_memory[12061] = 3'b000;
        rom_memory[12062] = 3'b000;
        rom_memory[12063] = 3'b000;
        rom_memory[12064] = 3'b000;
        rom_memory[12065] = 3'b000;
        rom_memory[12066] = 3'b000;
        rom_memory[12067] = 3'b000;
        rom_memory[12068] = 3'b000;
        rom_memory[12069] = 3'b000;
        rom_memory[12070] = 3'b000;
        rom_memory[12071] = 3'b000;
        rom_memory[12072] = 3'b000;
        rom_memory[12073] = 3'b000;
        rom_memory[12074] = 3'b000;
        rom_memory[12075] = 3'b000;
        rom_memory[12076] = 3'b000;
        rom_memory[12077] = 3'b000;
        rom_memory[12078] = 3'b000;
        rom_memory[12079] = 3'b000;
        rom_memory[12080] = 3'b000;
        rom_memory[12081] = 3'b010;
        rom_memory[12082] = 3'b000;
        rom_memory[12083] = 3'b000;
        rom_memory[12084] = 3'b000;
        rom_memory[12085] = 3'b010;
        rom_memory[12086] = 3'b000;
        rom_memory[12087] = 3'b000;
        rom_memory[12088] = 3'b011;
        rom_memory[12089] = 3'b011;
        rom_memory[12090] = 3'b011;
        rom_memory[12091] = 3'b011;
        rom_memory[12092] = 3'b011;
        rom_memory[12093] = 3'b011;
        rom_memory[12094] = 3'b011;
        rom_memory[12095] = 3'b011;
        rom_memory[12096] = 3'b011;
        rom_memory[12097] = 3'b011;
        rom_memory[12098] = 3'b011;
        rom_memory[12099] = 3'b011;
        rom_memory[12100] = 3'b001;
        rom_memory[12101] = 3'b001;
        rom_memory[12102] = 3'b111;
        rom_memory[12103] = 3'b111;
        rom_memory[12104] = 3'b110;
        rom_memory[12105] = 3'b110;
        rom_memory[12106] = 3'b110;
        rom_memory[12107] = 3'b110;
        rom_memory[12108] = 3'b110;
        rom_memory[12109] = 3'b110;
        rom_memory[12110] = 3'b110;
        rom_memory[12111] = 3'b110;
        rom_memory[12112] = 3'b110;
        rom_memory[12113] = 3'b110;
        rom_memory[12114] = 3'b110;
        rom_memory[12115] = 3'b110;
        rom_memory[12116] = 3'b110;
        rom_memory[12117] = 3'b110;
        rom_memory[12118] = 3'b110;
        rom_memory[12119] = 3'b110;
        rom_memory[12120] = 3'b110;
        rom_memory[12121] = 3'b110;
        rom_memory[12122] = 3'b110;
        rom_memory[12123] = 3'b110;
        rom_memory[12124] = 3'b110;
        rom_memory[12125] = 3'b110;
        rom_memory[12126] = 3'b110;
        rom_memory[12127] = 3'b110;
        rom_memory[12128] = 3'b110;
        rom_memory[12129] = 3'b110;
        rom_memory[12130] = 3'b110;
        rom_memory[12131] = 3'b110;
        rom_memory[12132] = 3'b110;
        rom_memory[12133] = 3'b110;
        rom_memory[12134] = 3'b110;
        rom_memory[12135] = 3'b110;
        rom_memory[12136] = 3'b110;
        rom_memory[12137] = 3'b110;
        rom_memory[12138] = 3'b110;
        rom_memory[12139] = 3'b110;
        rom_memory[12140] = 3'b110;
        rom_memory[12141] = 3'b110;
        rom_memory[12142] = 3'b110;
        rom_memory[12143] = 3'b110;
        rom_memory[12144] = 3'b110;
        rom_memory[12145] = 3'b110;
        rom_memory[12146] = 3'b110;
        rom_memory[12147] = 3'b110;
        rom_memory[12148] = 3'b110;
        rom_memory[12149] = 3'b110;
        rom_memory[12150] = 3'b110;
        rom_memory[12151] = 3'b110;
        rom_memory[12152] = 3'b110;
        rom_memory[12153] = 3'b110;
        rom_memory[12154] = 3'b110;
        rom_memory[12155] = 3'b110;
        rom_memory[12156] = 3'b110;
        rom_memory[12157] = 3'b110;
        rom_memory[12158] = 3'b110;
        rom_memory[12159] = 3'b110;
        rom_memory[12160] = 3'b110;
        rom_memory[12161] = 3'b110;
        rom_memory[12162] = 3'b110;
        rom_memory[12163] = 3'b110;
        rom_memory[12164] = 3'b110;
        rom_memory[12165] = 3'b110;
        rom_memory[12166] = 3'b110;
        rom_memory[12167] = 3'b110;
        rom_memory[12168] = 3'b110;
        rom_memory[12169] = 3'b110;
        rom_memory[12170] = 3'b110;
        rom_memory[12171] = 3'b110;
        rom_memory[12172] = 3'b110;
        rom_memory[12173] = 3'b110;
        rom_memory[12174] = 3'b110;
        rom_memory[12175] = 3'b110;
        rom_memory[12176] = 3'b110;
        rom_memory[12177] = 3'b110;
        rom_memory[12178] = 3'b110;
        rom_memory[12179] = 3'b110;
        rom_memory[12180] = 3'b110;
        rom_memory[12181] = 3'b110;
        rom_memory[12182] = 3'b110;
        rom_memory[12183] = 3'b110;
        rom_memory[12184] = 3'b110;
        rom_memory[12185] = 3'b110;
        rom_memory[12186] = 3'b110;
        rom_memory[12187] = 3'b110;
        rom_memory[12188] = 3'b110;
        rom_memory[12189] = 3'b110;
        rom_memory[12190] = 3'b110;
        rom_memory[12191] = 3'b110;
        rom_memory[12192] = 3'b110;
        rom_memory[12193] = 3'b110;
        rom_memory[12194] = 3'b110;
        rom_memory[12195] = 3'b110;
        rom_memory[12196] = 3'b110;
        rom_memory[12197] = 3'b110;
        rom_memory[12198] = 3'b110;
        rom_memory[12199] = 3'b110;
        rom_memory[12200] = 3'b110;
        rom_memory[12201] = 3'b110;
        rom_memory[12202] = 3'b110;
        rom_memory[12203] = 3'b110;
        rom_memory[12204] = 3'b110;
        rom_memory[12205] = 3'b110;
        rom_memory[12206] = 3'b110;
        rom_memory[12207] = 3'b110;
        rom_memory[12208] = 3'b110;
        rom_memory[12209] = 3'b110;
        rom_memory[12210] = 3'b110;
        rom_memory[12211] = 3'b110;
        rom_memory[12212] = 3'b110;
        rom_memory[12213] = 3'b110;
        rom_memory[12214] = 3'b110;
        rom_memory[12215] = 3'b110;
        rom_memory[12216] = 3'b110;
        rom_memory[12217] = 3'b110;
        rom_memory[12218] = 3'b110;
        rom_memory[12219] = 3'b110;
        rom_memory[12220] = 3'b110;
        rom_memory[12221] = 3'b110;
        rom_memory[12222] = 3'b110;
        rom_memory[12223] = 3'b110;
        rom_memory[12224] = 3'b110;
        rom_memory[12225] = 3'b110;
        rom_memory[12226] = 3'b110;
        rom_memory[12227] = 3'b110;
        rom_memory[12228] = 3'b110;
        rom_memory[12229] = 3'b110;
        rom_memory[12230] = 3'b110;
        rom_memory[12231] = 3'b110;
        rom_memory[12232] = 3'b110;
        rom_memory[12233] = 3'b110;
        rom_memory[12234] = 3'b110;
        rom_memory[12235] = 3'b110;
        rom_memory[12236] = 3'b110;
        rom_memory[12237] = 3'b110;
        rom_memory[12238] = 3'b110;
        rom_memory[12239] = 3'b110;
        rom_memory[12240] = 3'b110;
        rom_memory[12241] = 3'b110;
        rom_memory[12242] = 3'b110;
        rom_memory[12243] = 3'b110;
        rom_memory[12244] = 3'b110;
        rom_memory[12245] = 3'b110;
        rom_memory[12246] = 3'b110;
        rom_memory[12247] = 3'b110;
        rom_memory[12248] = 3'b110;
        rom_memory[12249] = 3'b110;
        rom_memory[12250] = 3'b110;
        rom_memory[12251] = 3'b110;
        rom_memory[12252] = 3'b110;
        rom_memory[12253] = 3'b110;
        rom_memory[12254] = 3'b110;
        rom_memory[12255] = 3'b110;
        rom_memory[12256] = 3'b110;
        rom_memory[12257] = 3'b110;
        rom_memory[12258] = 3'b110;
        rom_memory[12259] = 3'b110;
        rom_memory[12260] = 3'b110;
        rom_memory[12261] = 3'b110;
        rom_memory[12262] = 3'b110;
        rom_memory[12263] = 3'b110;
        rom_memory[12264] = 3'b110;
        rom_memory[12265] = 3'b110;
        rom_memory[12266] = 3'b110;
        rom_memory[12267] = 3'b110;
        rom_memory[12268] = 3'b110;
        rom_memory[12269] = 3'b110;
        rom_memory[12270] = 3'b110;
        rom_memory[12271] = 3'b110;
        rom_memory[12272] = 3'b110;
        rom_memory[12273] = 3'b110;
        rom_memory[12274] = 3'b110;
        rom_memory[12275] = 3'b110;
        rom_memory[12276] = 3'b110;
        rom_memory[12277] = 3'b110;
        rom_memory[12278] = 3'b110;
        rom_memory[12279] = 3'b110;
        rom_memory[12280] = 3'b110;
        rom_memory[12281] = 3'b110;
        rom_memory[12282] = 3'b111;
        rom_memory[12283] = 3'b110;
        rom_memory[12284] = 3'b111;
        rom_memory[12285] = 3'b111;
        rom_memory[12286] = 3'b111;
        rom_memory[12287] = 3'b111;
        rom_memory[12288] = 3'b000;
        rom_memory[12289] = 3'b000;
        rom_memory[12290] = 3'b000;
        rom_memory[12291] = 3'b000;
        rom_memory[12292] = 3'b000;
        rom_memory[12293] = 3'b000;
        rom_memory[12294] = 3'b000;
        rom_memory[12295] = 3'b000;
        rom_memory[12296] = 3'b000;
        rom_memory[12297] = 3'b000;
        rom_memory[12298] = 3'b000;
        rom_memory[12299] = 3'b000;
        rom_memory[12300] = 3'b000;
        rom_memory[12301] = 3'b000;
        rom_memory[12302] = 3'b000;
        rom_memory[12303] = 3'b000;
        rom_memory[12304] = 3'b000;
        rom_memory[12305] = 3'b000;
        rom_memory[12306] = 3'b000;
        rom_memory[12307] = 3'b000;
        rom_memory[12308] = 3'b000;
        rom_memory[12309] = 3'b000;
        rom_memory[12310] = 3'b000;
        rom_memory[12311] = 3'b000;
        rom_memory[12312] = 3'b000;
        rom_memory[12313] = 3'b000;
        rom_memory[12314] = 3'b000;
        rom_memory[12315] = 3'b000;
        rom_memory[12316] = 3'b000;
        rom_memory[12317] = 3'b000;
        rom_memory[12318] = 3'b000;
        rom_memory[12319] = 3'b000;
        rom_memory[12320] = 3'b000;
        rom_memory[12321] = 3'b000;
        rom_memory[12322] = 3'b000;
        rom_memory[12323] = 3'b000;
        rom_memory[12324] = 3'b000;
        rom_memory[12325] = 3'b000;
        rom_memory[12326] = 3'b000;
        rom_memory[12327] = 3'b000;
        rom_memory[12328] = 3'b000;
        rom_memory[12329] = 3'b000;
        rom_memory[12330] = 3'b011;
        rom_memory[12331] = 3'b011;
        rom_memory[12332] = 3'b011;
        rom_memory[12333] = 3'b011;
        rom_memory[12334] = 3'b011;
        rom_memory[12335] = 3'b001;
        rom_memory[12336] = 3'b011;
        rom_memory[12337] = 3'b011;
        rom_memory[12338] = 3'b011;
        rom_memory[12339] = 3'b011;
        rom_memory[12340] = 3'b011;
        rom_memory[12341] = 3'b001;
        rom_memory[12342] = 3'b111;
        rom_memory[12343] = 3'b111;
        rom_memory[12344] = 3'b110;
        rom_memory[12345] = 3'b110;
        rom_memory[12346] = 3'b110;
        rom_memory[12347] = 3'b110;
        rom_memory[12348] = 3'b110;
        rom_memory[12349] = 3'b110;
        rom_memory[12350] = 3'b110;
        rom_memory[12351] = 3'b110;
        rom_memory[12352] = 3'b110;
        rom_memory[12353] = 3'b110;
        rom_memory[12354] = 3'b110;
        rom_memory[12355] = 3'b110;
        rom_memory[12356] = 3'b110;
        rom_memory[12357] = 3'b110;
        rom_memory[12358] = 3'b110;
        rom_memory[12359] = 3'b110;
        rom_memory[12360] = 3'b110;
        rom_memory[12361] = 3'b110;
        rom_memory[12362] = 3'b110;
        rom_memory[12363] = 3'b110;
        rom_memory[12364] = 3'b110;
        rom_memory[12365] = 3'b110;
        rom_memory[12366] = 3'b110;
        rom_memory[12367] = 3'b110;
        rom_memory[12368] = 3'b110;
        rom_memory[12369] = 3'b110;
        rom_memory[12370] = 3'b110;
        rom_memory[12371] = 3'b110;
        rom_memory[12372] = 3'b110;
        rom_memory[12373] = 3'b110;
        rom_memory[12374] = 3'b110;
        rom_memory[12375] = 3'b110;
        rom_memory[12376] = 3'b110;
        rom_memory[12377] = 3'b111;
        rom_memory[12378] = 3'b110;
        rom_memory[12379] = 3'b110;
        rom_memory[12380] = 3'b110;
        rom_memory[12381] = 3'b110;
        rom_memory[12382] = 3'b110;
        rom_memory[12383] = 3'b111;
        rom_memory[12384] = 3'b110;
        rom_memory[12385] = 3'b110;
        rom_memory[12386] = 3'b110;
        rom_memory[12387] = 3'b110;
        rom_memory[12388] = 3'b110;
        rom_memory[12389] = 3'b110;
        rom_memory[12390] = 3'b110;
        rom_memory[12391] = 3'b110;
        rom_memory[12392] = 3'b110;
        rom_memory[12393] = 3'b110;
        rom_memory[12394] = 3'b110;
        rom_memory[12395] = 3'b110;
        rom_memory[12396] = 3'b110;
        rom_memory[12397] = 3'b110;
        rom_memory[12398] = 3'b110;
        rom_memory[12399] = 3'b110;
        rom_memory[12400] = 3'b110;
        rom_memory[12401] = 3'b110;
        rom_memory[12402] = 3'b110;
        rom_memory[12403] = 3'b110;
        rom_memory[12404] = 3'b110;
        rom_memory[12405] = 3'b110;
        rom_memory[12406] = 3'b110;
        rom_memory[12407] = 3'b110;
        rom_memory[12408] = 3'b110;
        rom_memory[12409] = 3'b110;
        rom_memory[12410] = 3'b110;
        rom_memory[12411] = 3'b110;
        rom_memory[12412] = 3'b110;
        rom_memory[12413] = 3'b110;
        rom_memory[12414] = 3'b110;
        rom_memory[12415] = 3'b110;
        rom_memory[12416] = 3'b110;
        rom_memory[12417] = 3'b110;
        rom_memory[12418] = 3'b110;
        rom_memory[12419] = 3'b110;
        rom_memory[12420] = 3'b110;
        rom_memory[12421] = 3'b110;
        rom_memory[12422] = 3'b110;
        rom_memory[12423] = 3'b110;
        rom_memory[12424] = 3'b110;
        rom_memory[12425] = 3'b110;
        rom_memory[12426] = 3'b110;
        rom_memory[12427] = 3'b110;
        rom_memory[12428] = 3'b110;
        rom_memory[12429] = 3'b110;
        rom_memory[12430] = 3'b110;
        rom_memory[12431] = 3'b110;
        rom_memory[12432] = 3'b110;
        rom_memory[12433] = 3'b110;
        rom_memory[12434] = 3'b110;
        rom_memory[12435] = 3'b110;
        rom_memory[12436] = 3'b110;
        rom_memory[12437] = 3'b110;
        rom_memory[12438] = 3'b110;
        rom_memory[12439] = 3'b110;
        rom_memory[12440] = 3'b110;
        rom_memory[12441] = 3'b110;
        rom_memory[12442] = 3'b110;
        rom_memory[12443] = 3'b110;
        rom_memory[12444] = 3'b110;
        rom_memory[12445] = 3'b110;
        rom_memory[12446] = 3'b110;
        rom_memory[12447] = 3'b110;
        rom_memory[12448] = 3'b110;
        rom_memory[12449] = 3'b110;
        rom_memory[12450] = 3'b110;
        rom_memory[12451] = 3'b110;
        rom_memory[12452] = 3'b110;
        rom_memory[12453] = 3'b110;
        rom_memory[12454] = 3'b110;
        rom_memory[12455] = 3'b110;
        rom_memory[12456] = 3'b110;
        rom_memory[12457] = 3'b110;
        rom_memory[12458] = 3'b110;
        rom_memory[12459] = 3'b110;
        rom_memory[12460] = 3'b110;
        rom_memory[12461] = 3'b110;
        rom_memory[12462] = 3'b110;
        rom_memory[12463] = 3'b110;
        rom_memory[12464] = 3'b110;
        rom_memory[12465] = 3'b110;
        rom_memory[12466] = 3'b110;
        rom_memory[12467] = 3'b110;
        rom_memory[12468] = 3'b110;
        rom_memory[12469] = 3'b110;
        rom_memory[12470] = 3'b110;
        rom_memory[12471] = 3'b110;
        rom_memory[12472] = 3'b110;
        rom_memory[12473] = 3'b110;
        rom_memory[12474] = 3'b110;
        rom_memory[12475] = 3'b110;
        rom_memory[12476] = 3'b110;
        rom_memory[12477] = 3'b110;
        rom_memory[12478] = 3'b110;
        rom_memory[12479] = 3'b110;
        rom_memory[12480] = 3'b110;
        rom_memory[12481] = 3'b110;
        rom_memory[12482] = 3'b110;
        rom_memory[12483] = 3'b110;
        rom_memory[12484] = 3'b110;
        rom_memory[12485] = 3'b110;
        rom_memory[12486] = 3'b110;
        rom_memory[12487] = 3'b110;
        rom_memory[12488] = 3'b110;
        rom_memory[12489] = 3'b110;
        rom_memory[12490] = 3'b110;
        rom_memory[12491] = 3'b110;
        rom_memory[12492] = 3'b110;
        rom_memory[12493] = 3'b110;
        rom_memory[12494] = 3'b110;
        rom_memory[12495] = 3'b110;
        rom_memory[12496] = 3'b110;
        rom_memory[12497] = 3'b110;
        rom_memory[12498] = 3'b110;
        rom_memory[12499] = 3'b110;
        rom_memory[12500] = 3'b110;
        rom_memory[12501] = 3'b110;
        rom_memory[12502] = 3'b110;
        rom_memory[12503] = 3'b110;
        rom_memory[12504] = 3'b110;
        rom_memory[12505] = 3'b110;
        rom_memory[12506] = 3'b110;
        rom_memory[12507] = 3'b110;
        rom_memory[12508] = 3'b110;
        rom_memory[12509] = 3'b110;
        rom_memory[12510] = 3'b110;
        rom_memory[12511] = 3'b110;
        rom_memory[12512] = 3'b110;
        rom_memory[12513] = 3'b110;
        rom_memory[12514] = 3'b110;
        rom_memory[12515] = 3'b110;
        rom_memory[12516] = 3'b110;
        rom_memory[12517] = 3'b110;
        rom_memory[12518] = 3'b110;
        rom_memory[12519] = 3'b110;
        rom_memory[12520] = 3'b110;
        rom_memory[12521] = 3'b110;
        rom_memory[12522] = 3'b111;
        rom_memory[12523] = 3'b111;
        rom_memory[12524] = 3'b111;
        rom_memory[12525] = 3'b111;
        rom_memory[12526] = 3'b111;
        rom_memory[12527] = 3'b111;
        rom_memory[12528] = 3'b111;
        rom_memory[12529] = 3'b000;
        rom_memory[12530] = 3'b000;
        rom_memory[12531] = 3'b000;
        rom_memory[12532] = 3'b000;
        rom_memory[12533] = 3'b000;
        rom_memory[12534] = 3'b000;
        rom_memory[12535] = 3'b000;
        rom_memory[12536] = 3'b000;
        rom_memory[12537] = 3'b000;
        rom_memory[12538] = 3'b000;
        rom_memory[12539] = 3'b000;
        rom_memory[12540] = 3'b000;
        rom_memory[12541] = 3'b000;
        rom_memory[12542] = 3'b000;
        rom_memory[12543] = 3'b000;
        rom_memory[12544] = 3'b000;
        rom_memory[12545] = 3'b000;
        rom_memory[12546] = 3'b000;
        rom_memory[12547] = 3'b000;
        rom_memory[12548] = 3'b000;
        rom_memory[12549] = 3'b000;
        rom_memory[12550] = 3'b000;
        rom_memory[12551] = 3'b000;
        rom_memory[12552] = 3'b000;
        rom_memory[12553] = 3'b000;
        rom_memory[12554] = 3'b000;
        rom_memory[12555] = 3'b000;
        rom_memory[12556] = 3'b000;
        rom_memory[12557] = 3'b000;
        rom_memory[12558] = 3'b000;
        rom_memory[12559] = 3'b000;
        rom_memory[12560] = 3'b000;
        rom_memory[12561] = 3'b000;
        rom_memory[12562] = 3'b000;
        rom_memory[12563] = 3'b000;
        rom_memory[12564] = 3'b000;
        rom_memory[12565] = 3'b000;
        rom_memory[12566] = 3'b011;
        rom_memory[12567] = 3'b000;
        rom_memory[12568] = 3'b000;
        rom_memory[12569] = 3'b000;
        rom_memory[12570] = 3'b011;
        rom_memory[12571] = 3'b011;
        rom_memory[12572] = 3'b011;
        rom_memory[12573] = 3'b011;
        rom_memory[12574] = 3'b011;
        rom_memory[12575] = 3'b011;
        rom_memory[12576] = 3'b011;
        rom_memory[12577] = 3'b011;
        rom_memory[12578] = 3'b011;
        rom_memory[12579] = 3'b011;
        rom_memory[12580] = 3'b011;
        rom_memory[12581] = 3'b011;
        rom_memory[12582] = 3'b011;
        rom_memory[12583] = 3'b111;
        rom_memory[12584] = 3'b111;
        rom_memory[12585] = 3'b110;
        rom_memory[12586] = 3'b110;
        rom_memory[12587] = 3'b110;
        rom_memory[12588] = 3'b110;
        rom_memory[12589] = 3'b110;
        rom_memory[12590] = 3'b110;
        rom_memory[12591] = 3'b110;
        rom_memory[12592] = 3'b110;
        rom_memory[12593] = 3'b110;
        rom_memory[12594] = 3'b110;
        rom_memory[12595] = 3'b110;
        rom_memory[12596] = 3'b110;
        rom_memory[12597] = 3'b110;
        rom_memory[12598] = 3'b110;
        rom_memory[12599] = 3'b110;
        rom_memory[12600] = 3'b110;
        rom_memory[12601] = 3'b110;
        rom_memory[12602] = 3'b110;
        rom_memory[12603] = 3'b110;
        rom_memory[12604] = 3'b110;
        rom_memory[12605] = 3'b111;
        rom_memory[12606] = 3'b110;
        rom_memory[12607] = 3'b110;
        rom_memory[12608] = 3'b110;
        rom_memory[12609] = 3'b110;
        rom_memory[12610] = 3'b110;
        rom_memory[12611] = 3'b110;
        rom_memory[12612] = 3'b110;
        rom_memory[12613] = 3'b110;
        rom_memory[12614] = 3'b110;
        rom_memory[12615] = 3'b110;
        rom_memory[12616] = 3'b111;
        rom_memory[12617] = 3'b111;
        rom_memory[12618] = 3'b110;
        rom_memory[12619] = 3'b110;
        rom_memory[12620] = 3'b110;
        rom_memory[12621] = 3'b110;
        rom_memory[12622] = 3'b110;
        rom_memory[12623] = 3'b110;
        rom_memory[12624] = 3'b110;
        rom_memory[12625] = 3'b110;
        rom_memory[12626] = 3'b110;
        rom_memory[12627] = 3'b110;
        rom_memory[12628] = 3'b110;
        rom_memory[12629] = 3'b110;
        rom_memory[12630] = 3'b110;
        rom_memory[12631] = 3'b110;
        rom_memory[12632] = 3'b110;
        rom_memory[12633] = 3'b110;
        rom_memory[12634] = 3'b110;
        rom_memory[12635] = 3'b110;
        rom_memory[12636] = 3'b110;
        rom_memory[12637] = 3'b110;
        rom_memory[12638] = 3'b110;
        rom_memory[12639] = 3'b110;
        rom_memory[12640] = 3'b110;
        rom_memory[12641] = 3'b110;
        rom_memory[12642] = 3'b110;
        rom_memory[12643] = 3'b110;
        rom_memory[12644] = 3'b110;
        rom_memory[12645] = 3'b110;
        rom_memory[12646] = 3'b110;
        rom_memory[12647] = 3'b110;
        rom_memory[12648] = 3'b110;
        rom_memory[12649] = 3'b110;
        rom_memory[12650] = 3'b110;
        rom_memory[12651] = 3'b110;
        rom_memory[12652] = 3'b110;
        rom_memory[12653] = 3'b110;
        rom_memory[12654] = 3'b110;
        rom_memory[12655] = 3'b110;
        rom_memory[12656] = 3'b110;
        rom_memory[12657] = 3'b110;
        rom_memory[12658] = 3'b110;
        rom_memory[12659] = 3'b110;
        rom_memory[12660] = 3'b110;
        rom_memory[12661] = 3'b110;
        rom_memory[12662] = 3'b110;
        rom_memory[12663] = 3'b110;
        rom_memory[12664] = 3'b110;
        rom_memory[12665] = 3'b110;
        rom_memory[12666] = 3'b110;
        rom_memory[12667] = 3'b110;
        rom_memory[12668] = 3'b110;
        rom_memory[12669] = 3'b110;
        rom_memory[12670] = 3'b110;
        rom_memory[12671] = 3'b110;
        rom_memory[12672] = 3'b110;
        rom_memory[12673] = 3'b110;
        rom_memory[12674] = 3'b110;
        rom_memory[12675] = 3'b110;
        rom_memory[12676] = 3'b110;
        rom_memory[12677] = 3'b110;
        rom_memory[12678] = 3'b110;
        rom_memory[12679] = 3'b110;
        rom_memory[12680] = 3'b110;
        rom_memory[12681] = 3'b110;
        rom_memory[12682] = 3'b110;
        rom_memory[12683] = 3'b110;
        rom_memory[12684] = 3'b110;
        rom_memory[12685] = 3'b110;
        rom_memory[12686] = 3'b110;
        rom_memory[12687] = 3'b110;
        rom_memory[12688] = 3'b110;
        rom_memory[12689] = 3'b110;
        rom_memory[12690] = 3'b110;
        rom_memory[12691] = 3'b110;
        rom_memory[12692] = 3'b110;
        rom_memory[12693] = 3'b110;
        rom_memory[12694] = 3'b110;
        rom_memory[12695] = 3'b110;
        rom_memory[12696] = 3'b110;
        rom_memory[12697] = 3'b110;
        rom_memory[12698] = 3'b110;
        rom_memory[12699] = 3'b110;
        rom_memory[12700] = 3'b110;
        rom_memory[12701] = 3'b110;
        rom_memory[12702] = 3'b110;
        rom_memory[12703] = 3'b110;
        rom_memory[12704] = 3'b110;
        rom_memory[12705] = 3'b110;
        rom_memory[12706] = 3'b110;
        rom_memory[12707] = 3'b110;
        rom_memory[12708] = 3'b110;
        rom_memory[12709] = 3'b110;
        rom_memory[12710] = 3'b110;
        rom_memory[12711] = 3'b110;
        rom_memory[12712] = 3'b110;
        rom_memory[12713] = 3'b110;
        rom_memory[12714] = 3'b110;
        rom_memory[12715] = 3'b110;
        rom_memory[12716] = 3'b110;
        rom_memory[12717] = 3'b110;
        rom_memory[12718] = 3'b110;
        rom_memory[12719] = 3'b110;
        rom_memory[12720] = 3'b110;
        rom_memory[12721] = 3'b110;
        rom_memory[12722] = 3'b110;
        rom_memory[12723] = 3'b110;
        rom_memory[12724] = 3'b110;
        rom_memory[12725] = 3'b110;
        rom_memory[12726] = 3'b110;
        rom_memory[12727] = 3'b110;
        rom_memory[12728] = 3'b110;
        rom_memory[12729] = 3'b110;
        rom_memory[12730] = 3'b110;
        rom_memory[12731] = 3'b110;
        rom_memory[12732] = 3'b110;
        rom_memory[12733] = 3'b110;
        rom_memory[12734] = 3'b110;
        rom_memory[12735] = 3'b110;
        rom_memory[12736] = 3'b110;
        rom_memory[12737] = 3'b110;
        rom_memory[12738] = 3'b110;
        rom_memory[12739] = 3'b110;
        rom_memory[12740] = 3'b110;
        rom_memory[12741] = 3'b110;
        rom_memory[12742] = 3'b110;
        rom_memory[12743] = 3'b110;
        rom_memory[12744] = 3'b110;
        rom_memory[12745] = 3'b110;
        rom_memory[12746] = 3'b110;
        rom_memory[12747] = 3'b110;
        rom_memory[12748] = 3'b110;
        rom_memory[12749] = 3'b110;
        rom_memory[12750] = 3'b110;
        rom_memory[12751] = 3'b110;
        rom_memory[12752] = 3'b110;
        rom_memory[12753] = 3'b110;
        rom_memory[12754] = 3'b110;
        rom_memory[12755] = 3'b110;
        rom_memory[12756] = 3'b110;
        rom_memory[12757] = 3'b110;
        rom_memory[12758] = 3'b110;
        rom_memory[12759] = 3'b110;
        rom_memory[12760] = 3'b110;
        rom_memory[12761] = 3'b111;
        rom_memory[12762] = 3'b111;
        rom_memory[12763] = 3'b111;
        rom_memory[12764] = 3'b111;
        rom_memory[12765] = 3'b111;
        rom_memory[12766] = 3'b111;
        rom_memory[12767] = 3'b111;
        rom_memory[12768] = 3'b111;
        rom_memory[12769] = 3'b000;
        rom_memory[12770] = 3'b000;
        rom_memory[12771] = 3'b000;
        rom_memory[12772] = 3'b000;
        rom_memory[12773] = 3'b000;
        rom_memory[12774] = 3'b000;
        rom_memory[12775] = 3'b000;
        rom_memory[12776] = 3'b000;
        rom_memory[12777] = 3'b000;
        rom_memory[12778] = 3'b000;
        rom_memory[12779] = 3'b000;
        rom_memory[12780] = 3'b000;
        rom_memory[12781] = 3'b000;
        rom_memory[12782] = 3'b000;
        rom_memory[12783] = 3'b000;
        rom_memory[12784] = 3'b000;
        rom_memory[12785] = 3'b000;
        rom_memory[12786] = 3'b000;
        rom_memory[12787] = 3'b000;
        rom_memory[12788] = 3'b000;
        rom_memory[12789] = 3'b000;
        rom_memory[12790] = 3'b000;
        rom_memory[12791] = 3'b000;
        rom_memory[12792] = 3'b000;
        rom_memory[12793] = 3'b000;
        rom_memory[12794] = 3'b000;
        rom_memory[12795] = 3'b000;
        rom_memory[12796] = 3'b000;
        rom_memory[12797] = 3'b011;
        rom_memory[12798] = 3'b000;
        rom_memory[12799] = 3'b000;
        rom_memory[12800] = 3'b000;
        rom_memory[12801] = 3'b000;
        rom_memory[12802] = 3'b000;
        rom_memory[12803] = 3'b011;
        rom_memory[12804] = 3'b011;
        rom_memory[12805] = 3'b000;
        rom_memory[12806] = 3'b010;
        rom_memory[12807] = 3'b000;
        rom_memory[12808] = 3'b010;
        rom_memory[12809] = 3'b011;
        rom_memory[12810] = 3'b111;
        rom_memory[12811] = 3'b111;
        rom_memory[12812] = 3'b111;
        rom_memory[12813] = 3'b111;
        rom_memory[12814] = 3'b011;
        rom_memory[12815] = 3'b011;
        rom_memory[12816] = 3'b011;
        rom_memory[12817] = 3'b011;
        rom_memory[12818] = 3'b011;
        rom_memory[12819] = 3'b011;
        rom_memory[12820] = 3'b011;
        rom_memory[12821] = 3'b001;
        rom_memory[12822] = 3'b001;
        rom_memory[12823] = 3'b111;
        rom_memory[12824] = 3'b111;
        rom_memory[12825] = 3'b111;
        rom_memory[12826] = 3'b110;
        rom_memory[12827] = 3'b110;
        rom_memory[12828] = 3'b110;
        rom_memory[12829] = 3'b110;
        rom_memory[12830] = 3'b110;
        rom_memory[12831] = 3'b110;
        rom_memory[12832] = 3'b110;
        rom_memory[12833] = 3'b110;
        rom_memory[12834] = 3'b110;
        rom_memory[12835] = 3'b110;
        rom_memory[12836] = 3'b110;
        rom_memory[12837] = 3'b110;
        rom_memory[12838] = 3'b110;
        rom_memory[12839] = 3'b110;
        rom_memory[12840] = 3'b110;
        rom_memory[12841] = 3'b110;
        rom_memory[12842] = 3'b110;
        rom_memory[12843] = 3'b110;
        rom_memory[12844] = 3'b110;
        rom_memory[12845] = 3'b110;
        rom_memory[12846] = 3'b110;
        rom_memory[12847] = 3'b110;
        rom_memory[12848] = 3'b110;
        rom_memory[12849] = 3'b110;
        rom_memory[12850] = 3'b110;
        rom_memory[12851] = 3'b110;
        rom_memory[12852] = 3'b111;
        rom_memory[12853] = 3'b110;
        rom_memory[12854] = 3'b110;
        rom_memory[12855] = 3'b110;
        rom_memory[12856] = 3'b111;
        rom_memory[12857] = 3'b110;
        rom_memory[12858] = 3'b111;
        rom_memory[12859] = 3'b111;
        rom_memory[12860] = 3'b111;
        rom_memory[12861] = 3'b110;
        rom_memory[12862] = 3'b110;
        rom_memory[12863] = 3'b110;
        rom_memory[12864] = 3'b110;
        rom_memory[12865] = 3'b110;
        rom_memory[12866] = 3'b110;
        rom_memory[12867] = 3'b110;
        rom_memory[12868] = 3'b110;
        rom_memory[12869] = 3'b110;
        rom_memory[12870] = 3'b110;
        rom_memory[12871] = 3'b110;
        rom_memory[12872] = 3'b110;
        rom_memory[12873] = 3'b110;
        rom_memory[12874] = 3'b110;
        rom_memory[12875] = 3'b110;
        rom_memory[12876] = 3'b110;
        rom_memory[12877] = 3'b110;
        rom_memory[12878] = 3'b110;
        rom_memory[12879] = 3'b110;
        rom_memory[12880] = 3'b110;
        rom_memory[12881] = 3'b110;
        rom_memory[12882] = 3'b110;
        rom_memory[12883] = 3'b110;
        rom_memory[12884] = 3'b110;
        rom_memory[12885] = 3'b110;
        rom_memory[12886] = 3'b110;
        rom_memory[12887] = 3'b110;
        rom_memory[12888] = 3'b110;
        rom_memory[12889] = 3'b110;
        rom_memory[12890] = 3'b110;
        rom_memory[12891] = 3'b110;
        rom_memory[12892] = 3'b110;
        rom_memory[12893] = 3'b110;
        rom_memory[12894] = 3'b110;
        rom_memory[12895] = 3'b110;
        rom_memory[12896] = 3'b110;
        rom_memory[12897] = 3'b110;
        rom_memory[12898] = 3'b110;
        rom_memory[12899] = 3'b110;
        rom_memory[12900] = 3'b110;
        rom_memory[12901] = 3'b110;
        rom_memory[12902] = 3'b110;
        rom_memory[12903] = 3'b110;
        rom_memory[12904] = 3'b110;
        rom_memory[12905] = 3'b110;
        rom_memory[12906] = 3'b110;
        rom_memory[12907] = 3'b110;
        rom_memory[12908] = 3'b110;
        rom_memory[12909] = 3'b110;
        rom_memory[12910] = 3'b110;
        rom_memory[12911] = 3'b110;
        rom_memory[12912] = 3'b110;
        rom_memory[12913] = 3'b110;
        rom_memory[12914] = 3'b110;
        rom_memory[12915] = 3'b110;
        rom_memory[12916] = 3'b110;
        rom_memory[12917] = 3'b110;
        rom_memory[12918] = 3'b110;
        rom_memory[12919] = 3'b110;
        rom_memory[12920] = 3'b110;
        rom_memory[12921] = 3'b110;
        rom_memory[12922] = 3'b110;
        rom_memory[12923] = 3'b110;
        rom_memory[12924] = 3'b110;
        rom_memory[12925] = 3'b110;
        rom_memory[12926] = 3'b110;
        rom_memory[12927] = 3'b110;
        rom_memory[12928] = 3'b110;
        rom_memory[12929] = 3'b110;
        rom_memory[12930] = 3'b110;
        rom_memory[12931] = 3'b110;
        rom_memory[12932] = 3'b110;
        rom_memory[12933] = 3'b110;
        rom_memory[12934] = 3'b110;
        rom_memory[12935] = 3'b110;
        rom_memory[12936] = 3'b110;
        rom_memory[12937] = 3'b110;
        rom_memory[12938] = 3'b110;
        rom_memory[12939] = 3'b110;
        rom_memory[12940] = 3'b110;
        rom_memory[12941] = 3'b110;
        rom_memory[12942] = 3'b110;
        rom_memory[12943] = 3'b110;
        rom_memory[12944] = 3'b110;
        rom_memory[12945] = 3'b110;
        rom_memory[12946] = 3'b110;
        rom_memory[12947] = 3'b110;
        rom_memory[12948] = 3'b110;
        rom_memory[12949] = 3'b110;
        rom_memory[12950] = 3'b110;
        rom_memory[12951] = 3'b110;
        rom_memory[12952] = 3'b110;
        rom_memory[12953] = 3'b110;
        rom_memory[12954] = 3'b110;
        rom_memory[12955] = 3'b110;
        rom_memory[12956] = 3'b110;
        rom_memory[12957] = 3'b110;
        rom_memory[12958] = 3'b110;
        rom_memory[12959] = 3'b110;
        rom_memory[12960] = 3'b110;
        rom_memory[12961] = 3'b110;
        rom_memory[12962] = 3'b110;
        rom_memory[12963] = 3'b110;
        rom_memory[12964] = 3'b110;
        rom_memory[12965] = 3'b110;
        rom_memory[12966] = 3'b110;
        rom_memory[12967] = 3'b110;
        rom_memory[12968] = 3'b110;
        rom_memory[12969] = 3'b110;
        rom_memory[12970] = 3'b110;
        rom_memory[12971] = 3'b110;
        rom_memory[12972] = 3'b110;
        rom_memory[12973] = 3'b110;
        rom_memory[12974] = 3'b110;
        rom_memory[12975] = 3'b110;
        rom_memory[12976] = 3'b110;
        rom_memory[12977] = 3'b110;
        rom_memory[12978] = 3'b110;
        rom_memory[12979] = 3'b110;
        rom_memory[12980] = 3'b110;
        rom_memory[12981] = 3'b110;
        rom_memory[12982] = 3'b110;
        rom_memory[12983] = 3'b110;
        rom_memory[12984] = 3'b110;
        rom_memory[12985] = 3'b110;
        rom_memory[12986] = 3'b110;
        rom_memory[12987] = 3'b110;
        rom_memory[12988] = 3'b110;
        rom_memory[12989] = 3'b110;
        rom_memory[12990] = 3'b110;
        rom_memory[12991] = 3'b110;
        rom_memory[12992] = 3'b110;
        rom_memory[12993] = 3'b110;
        rom_memory[12994] = 3'b110;
        rom_memory[12995] = 3'b110;
        rom_memory[12996] = 3'b110;
        rom_memory[12997] = 3'b110;
        rom_memory[12998] = 3'b110;
        rom_memory[12999] = 3'b110;
        rom_memory[13000] = 3'b111;
        rom_memory[13001] = 3'b111;
        rom_memory[13002] = 3'b111;
        rom_memory[13003] = 3'b111;
        rom_memory[13004] = 3'b111;
        rom_memory[13005] = 3'b111;
        rom_memory[13006] = 3'b111;
        rom_memory[13007] = 3'b111;
        rom_memory[13008] = 3'b000;
        rom_memory[13009] = 3'b000;
        rom_memory[13010] = 3'b000;
        rom_memory[13011] = 3'b000;
        rom_memory[13012] = 3'b000;
        rom_memory[13013] = 3'b000;
        rom_memory[13014] = 3'b000;
        rom_memory[13015] = 3'b000;
        rom_memory[13016] = 3'b000;
        rom_memory[13017] = 3'b000;
        rom_memory[13018] = 3'b000;
        rom_memory[13019] = 3'b000;
        rom_memory[13020] = 3'b000;
        rom_memory[13021] = 3'b000;
        rom_memory[13022] = 3'b000;
        rom_memory[13023] = 3'b000;
        rom_memory[13024] = 3'b000;
        rom_memory[13025] = 3'b000;
        rom_memory[13026] = 3'b000;
        rom_memory[13027] = 3'b000;
        rom_memory[13028] = 3'b000;
        rom_memory[13029] = 3'b000;
        rom_memory[13030] = 3'b000;
        rom_memory[13031] = 3'b000;
        rom_memory[13032] = 3'b000;
        rom_memory[13033] = 3'b000;
        rom_memory[13034] = 3'b000;
        rom_memory[13035] = 3'b000;
        rom_memory[13036] = 3'b000;
        rom_memory[13037] = 3'b000;
        rom_memory[13038] = 3'b000;
        rom_memory[13039] = 3'b001;
        rom_memory[13040] = 3'b000;
        rom_memory[13041] = 3'b000;
        rom_memory[13042] = 3'b000;
        rom_memory[13043] = 3'b000;
        rom_memory[13044] = 3'b000;
        rom_memory[13045] = 3'b000;
        rom_memory[13046] = 3'b001;
        rom_memory[13047] = 3'b011;
        rom_memory[13048] = 3'b011;
        rom_memory[13049] = 3'b011;
        rom_memory[13050] = 3'b111;
        rom_memory[13051] = 3'b111;
        rom_memory[13052] = 3'b111;
        rom_memory[13053] = 3'b111;
        rom_memory[13054] = 3'b111;
        rom_memory[13055] = 3'b111;
        rom_memory[13056] = 3'b111;
        rom_memory[13057] = 3'b111;
        rom_memory[13058] = 3'b111;
        rom_memory[13059] = 3'b011;
        rom_memory[13060] = 3'b011;
        rom_memory[13061] = 3'b011;
        rom_memory[13062] = 3'b011;
        rom_memory[13063] = 3'b111;
        rom_memory[13064] = 3'b111;
        rom_memory[13065] = 3'b111;
        rom_memory[13066] = 3'b110;
        rom_memory[13067] = 3'b110;
        rom_memory[13068] = 3'b110;
        rom_memory[13069] = 3'b110;
        rom_memory[13070] = 3'b110;
        rom_memory[13071] = 3'b110;
        rom_memory[13072] = 3'b110;
        rom_memory[13073] = 3'b110;
        rom_memory[13074] = 3'b110;
        rom_memory[13075] = 3'b110;
        rom_memory[13076] = 3'b110;
        rom_memory[13077] = 3'b110;
        rom_memory[13078] = 3'b110;
        rom_memory[13079] = 3'b110;
        rom_memory[13080] = 3'b110;
        rom_memory[13081] = 3'b110;
        rom_memory[13082] = 3'b110;
        rom_memory[13083] = 3'b110;
        rom_memory[13084] = 3'b110;
        rom_memory[13085] = 3'b110;
        rom_memory[13086] = 3'b110;
        rom_memory[13087] = 3'b110;
        rom_memory[13088] = 3'b110;
        rom_memory[13089] = 3'b111;
        rom_memory[13090] = 3'b111;
        rom_memory[13091] = 3'b111;
        rom_memory[13092] = 3'b110;
        rom_memory[13093] = 3'b111;
        rom_memory[13094] = 3'b111;
        rom_memory[13095] = 3'b110;
        rom_memory[13096] = 3'b110;
        rom_memory[13097] = 3'b110;
        rom_memory[13098] = 3'b111;
        rom_memory[13099] = 3'b111;
        rom_memory[13100] = 3'b111;
        rom_memory[13101] = 3'b110;
        rom_memory[13102] = 3'b110;
        rom_memory[13103] = 3'b110;
        rom_memory[13104] = 3'b110;
        rom_memory[13105] = 3'b110;
        rom_memory[13106] = 3'b110;
        rom_memory[13107] = 3'b110;
        rom_memory[13108] = 3'b111;
        rom_memory[13109] = 3'b111;
        rom_memory[13110] = 3'b111;
        rom_memory[13111] = 3'b110;
        rom_memory[13112] = 3'b110;
        rom_memory[13113] = 3'b110;
        rom_memory[13114] = 3'b110;
        rom_memory[13115] = 3'b110;
        rom_memory[13116] = 3'b110;
        rom_memory[13117] = 3'b110;
        rom_memory[13118] = 3'b110;
        rom_memory[13119] = 3'b110;
        rom_memory[13120] = 3'b110;
        rom_memory[13121] = 3'b110;
        rom_memory[13122] = 3'b110;
        rom_memory[13123] = 3'b110;
        rom_memory[13124] = 3'b110;
        rom_memory[13125] = 3'b110;
        rom_memory[13126] = 3'b110;
        rom_memory[13127] = 3'b110;
        rom_memory[13128] = 3'b110;
        rom_memory[13129] = 3'b110;
        rom_memory[13130] = 3'b110;
        rom_memory[13131] = 3'b110;
        rom_memory[13132] = 3'b110;
        rom_memory[13133] = 3'b110;
        rom_memory[13134] = 3'b110;
        rom_memory[13135] = 3'b110;
        rom_memory[13136] = 3'b110;
        rom_memory[13137] = 3'b110;
        rom_memory[13138] = 3'b110;
        rom_memory[13139] = 3'b110;
        rom_memory[13140] = 3'b110;
        rom_memory[13141] = 3'b110;
        rom_memory[13142] = 3'b110;
        rom_memory[13143] = 3'b110;
        rom_memory[13144] = 3'b110;
        rom_memory[13145] = 3'b110;
        rom_memory[13146] = 3'b110;
        rom_memory[13147] = 3'b110;
        rom_memory[13148] = 3'b110;
        rom_memory[13149] = 3'b110;
        rom_memory[13150] = 3'b110;
        rom_memory[13151] = 3'b110;
        rom_memory[13152] = 3'b110;
        rom_memory[13153] = 3'b110;
        rom_memory[13154] = 3'b110;
        rom_memory[13155] = 3'b110;
        rom_memory[13156] = 3'b110;
        rom_memory[13157] = 3'b110;
        rom_memory[13158] = 3'b110;
        rom_memory[13159] = 3'b110;
        rom_memory[13160] = 3'b110;
        rom_memory[13161] = 3'b110;
        rom_memory[13162] = 3'b110;
        rom_memory[13163] = 3'b110;
        rom_memory[13164] = 3'b110;
        rom_memory[13165] = 3'b110;
        rom_memory[13166] = 3'b110;
        rom_memory[13167] = 3'b110;
        rom_memory[13168] = 3'b110;
        rom_memory[13169] = 3'b110;
        rom_memory[13170] = 3'b110;
        rom_memory[13171] = 3'b110;
        rom_memory[13172] = 3'b110;
        rom_memory[13173] = 3'b110;
        rom_memory[13174] = 3'b110;
        rom_memory[13175] = 3'b110;
        rom_memory[13176] = 3'b110;
        rom_memory[13177] = 3'b110;
        rom_memory[13178] = 3'b110;
        rom_memory[13179] = 3'b110;
        rom_memory[13180] = 3'b110;
        rom_memory[13181] = 3'b110;
        rom_memory[13182] = 3'b110;
        rom_memory[13183] = 3'b110;
        rom_memory[13184] = 3'b110;
        rom_memory[13185] = 3'b110;
        rom_memory[13186] = 3'b110;
        rom_memory[13187] = 3'b110;
        rom_memory[13188] = 3'b110;
        rom_memory[13189] = 3'b110;
        rom_memory[13190] = 3'b110;
        rom_memory[13191] = 3'b110;
        rom_memory[13192] = 3'b110;
        rom_memory[13193] = 3'b110;
        rom_memory[13194] = 3'b110;
        rom_memory[13195] = 3'b110;
        rom_memory[13196] = 3'b110;
        rom_memory[13197] = 3'b110;
        rom_memory[13198] = 3'b110;
        rom_memory[13199] = 3'b110;
        rom_memory[13200] = 3'b110;
        rom_memory[13201] = 3'b110;
        rom_memory[13202] = 3'b110;
        rom_memory[13203] = 3'b110;
        rom_memory[13204] = 3'b110;
        rom_memory[13205] = 3'b110;
        rom_memory[13206] = 3'b110;
        rom_memory[13207] = 3'b110;
        rom_memory[13208] = 3'b110;
        rom_memory[13209] = 3'b110;
        rom_memory[13210] = 3'b110;
        rom_memory[13211] = 3'b110;
        rom_memory[13212] = 3'b110;
        rom_memory[13213] = 3'b110;
        rom_memory[13214] = 3'b110;
        rom_memory[13215] = 3'b110;
        rom_memory[13216] = 3'b110;
        rom_memory[13217] = 3'b110;
        rom_memory[13218] = 3'b110;
        rom_memory[13219] = 3'b110;
        rom_memory[13220] = 3'b110;
        rom_memory[13221] = 3'b110;
        rom_memory[13222] = 3'b110;
        rom_memory[13223] = 3'b110;
        rom_memory[13224] = 3'b110;
        rom_memory[13225] = 3'b110;
        rom_memory[13226] = 3'b110;
        rom_memory[13227] = 3'b110;
        rom_memory[13228] = 3'b110;
        rom_memory[13229] = 3'b110;
        rom_memory[13230] = 3'b110;
        rom_memory[13231] = 3'b110;
        rom_memory[13232] = 3'b110;
        rom_memory[13233] = 3'b110;
        rom_memory[13234] = 3'b110;
        rom_memory[13235] = 3'b110;
        rom_memory[13236] = 3'b110;
        rom_memory[13237] = 3'b110;
        rom_memory[13238] = 3'b110;
        rom_memory[13239] = 3'b111;
        rom_memory[13240] = 3'b111;
        rom_memory[13241] = 3'b111;
        rom_memory[13242] = 3'b111;
        rom_memory[13243] = 3'b111;
        rom_memory[13244] = 3'b111;
        rom_memory[13245] = 3'b111;
        rom_memory[13246] = 3'b111;
        rom_memory[13247] = 3'b111;
        rom_memory[13248] = 3'b000;
        rom_memory[13249] = 3'b000;
        rom_memory[13250] = 3'b000;
        rom_memory[13251] = 3'b000;
        rom_memory[13252] = 3'b000;
        rom_memory[13253] = 3'b000;
        rom_memory[13254] = 3'b000;
        rom_memory[13255] = 3'b000;
        rom_memory[13256] = 3'b000;
        rom_memory[13257] = 3'b000;
        rom_memory[13258] = 3'b000;
        rom_memory[13259] = 3'b000;
        rom_memory[13260] = 3'b000;
        rom_memory[13261] = 3'b000;
        rom_memory[13262] = 3'b000;
        rom_memory[13263] = 3'b000;
        rom_memory[13264] = 3'b000;
        rom_memory[13265] = 3'b000;
        rom_memory[13266] = 3'b000;
        rom_memory[13267] = 3'b000;
        rom_memory[13268] = 3'b000;
        rom_memory[13269] = 3'b000;
        rom_memory[13270] = 3'b000;
        rom_memory[13271] = 3'b000;
        rom_memory[13272] = 3'b000;
        rom_memory[13273] = 3'b000;
        rom_memory[13274] = 3'b000;
        rom_memory[13275] = 3'b000;
        rom_memory[13276] = 3'b000;
        rom_memory[13277] = 3'b000;
        rom_memory[13278] = 3'b000;
        rom_memory[13279] = 3'b000;
        rom_memory[13280] = 3'b000;
        rom_memory[13281] = 3'b000;
        rom_memory[13282] = 3'b000;
        rom_memory[13283] = 3'b011;
        rom_memory[13284] = 3'b001;
        rom_memory[13285] = 3'b011;
        rom_memory[13286] = 3'b011;
        rom_memory[13287] = 3'b011;
        rom_memory[13288] = 3'b011;
        rom_memory[13289] = 3'b011;
        rom_memory[13290] = 3'b011;
        rom_memory[13291] = 3'b111;
        rom_memory[13292] = 3'b111;
        rom_memory[13293] = 3'b111;
        rom_memory[13294] = 3'b110;
        rom_memory[13295] = 3'b110;
        rom_memory[13296] = 3'b111;
        rom_memory[13297] = 3'b111;
        rom_memory[13298] = 3'b111;
        rom_memory[13299] = 3'b111;
        rom_memory[13300] = 3'b011;
        rom_memory[13301] = 3'b011;
        rom_memory[13302] = 3'b011;
        rom_memory[13303] = 3'b011;
        rom_memory[13304] = 3'b111;
        rom_memory[13305] = 3'b111;
        rom_memory[13306] = 3'b111;
        rom_memory[13307] = 3'b110;
        rom_memory[13308] = 3'b110;
        rom_memory[13309] = 3'b110;
        rom_memory[13310] = 3'b110;
        rom_memory[13311] = 3'b110;
        rom_memory[13312] = 3'b110;
        rom_memory[13313] = 3'b110;
        rom_memory[13314] = 3'b110;
        rom_memory[13315] = 3'b110;
        rom_memory[13316] = 3'b110;
        rom_memory[13317] = 3'b110;
        rom_memory[13318] = 3'b110;
        rom_memory[13319] = 3'b110;
        rom_memory[13320] = 3'b110;
        rom_memory[13321] = 3'b110;
        rom_memory[13322] = 3'b110;
        rom_memory[13323] = 3'b110;
        rom_memory[13324] = 3'b110;
        rom_memory[13325] = 3'b110;
        rom_memory[13326] = 3'b111;
        rom_memory[13327] = 3'b111;
        rom_memory[13328] = 3'b110;
        rom_memory[13329] = 3'b110;
        rom_memory[13330] = 3'b110;
        rom_memory[13331] = 3'b111;
        rom_memory[13332] = 3'b111;
        rom_memory[13333] = 3'b111;
        rom_memory[13334] = 3'b111;
        rom_memory[13335] = 3'b110;
        rom_memory[13336] = 3'b110;
        rom_memory[13337] = 3'b110;
        rom_memory[13338] = 3'b111;
        rom_memory[13339] = 3'b111;
        rom_memory[13340] = 3'b111;
        rom_memory[13341] = 3'b111;
        rom_memory[13342] = 3'b110;
        rom_memory[13343] = 3'b110;
        rom_memory[13344] = 3'b110;
        rom_memory[13345] = 3'b111;
        rom_memory[13346] = 3'b111;
        rom_memory[13347] = 3'b111;
        rom_memory[13348] = 3'b110;
        rom_memory[13349] = 3'b111;
        rom_memory[13350] = 3'b111;
        rom_memory[13351] = 3'b111;
        rom_memory[13352] = 3'b111;
        rom_memory[13353] = 3'b111;
        rom_memory[13354] = 3'b110;
        rom_memory[13355] = 3'b110;
        rom_memory[13356] = 3'b110;
        rom_memory[13357] = 3'b110;
        rom_memory[13358] = 3'b110;
        rom_memory[13359] = 3'b110;
        rom_memory[13360] = 3'b110;
        rom_memory[13361] = 3'b110;
        rom_memory[13362] = 3'b110;
        rom_memory[13363] = 3'b110;
        rom_memory[13364] = 3'b110;
        rom_memory[13365] = 3'b110;
        rom_memory[13366] = 3'b110;
        rom_memory[13367] = 3'b110;
        rom_memory[13368] = 3'b110;
        rom_memory[13369] = 3'b110;
        rom_memory[13370] = 3'b110;
        rom_memory[13371] = 3'b110;
        rom_memory[13372] = 3'b110;
        rom_memory[13373] = 3'b110;
        rom_memory[13374] = 3'b110;
        rom_memory[13375] = 3'b110;
        rom_memory[13376] = 3'b110;
        rom_memory[13377] = 3'b110;
        rom_memory[13378] = 3'b110;
        rom_memory[13379] = 3'b110;
        rom_memory[13380] = 3'b110;
        rom_memory[13381] = 3'b110;
        rom_memory[13382] = 3'b110;
        rom_memory[13383] = 3'b110;
        rom_memory[13384] = 3'b110;
        rom_memory[13385] = 3'b110;
        rom_memory[13386] = 3'b110;
        rom_memory[13387] = 3'b110;
        rom_memory[13388] = 3'b110;
        rom_memory[13389] = 3'b110;
        rom_memory[13390] = 3'b110;
        rom_memory[13391] = 3'b110;
        rom_memory[13392] = 3'b110;
        rom_memory[13393] = 3'b110;
        rom_memory[13394] = 3'b110;
        rom_memory[13395] = 3'b110;
        rom_memory[13396] = 3'b110;
        rom_memory[13397] = 3'b110;
        rom_memory[13398] = 3'b110;
        rom_memory[13399] = 3'b110;
        rom_memory[13400] = 3'b110;
        rom_memory[13401] = 3'b110;
        rom_memory[13402] = 3'b110;
        rom_memory[13403] = 3'b110;
        rom_memory[13404] = 3'b110;
        rom_memory[13405] = 3'b110;
        rom_memory[13406] = 3'b110;
        rom_memory[13407] = 3'b110;
        rom_memory[13408] = 3'b110;
        rom_memory[13409] = 3'b110;
        rom_memory[13410] = 3'b110;
        rom_memory[13411] = 3'b110;
        rom_memory[13412] = 3'b110;
        rom_memory[13413] = 3'b110;
        rom_memory[13414] = 3'b110;
        rom_memory[13415] = 3'b110;
        rom_memory[13416] = 3'b110;
        rom_memory[13417] = 3'b110;
        rom_memory[13418] = 3'b110;
        rom_memory[13419] = 3'b110;
        rom_memory[13420] = 3'b110;
        rom_memory[13421] = 3'b110;
        rom_memory[13422] = 3'b110;
        rom_memory[13423] = 3'b110;
        rom_memory[13424] = 3'b110;
        rom_memory[13425] = 3'b110;
        rom_memory[13426] = 3'b110;
        rom_memory[13427] = 3'b110;
        rom_memory[13428] = 3'b110;
        rom_memory[13429] = 3'b110;
        rom_memory[13430] = 3'b110;
        rom_memory[13431] = 3'b110;
        rom_memory[13432] = 3'b110;
        rom_memory[13433] = 3'b110;
        rom_memory[13434] = 3'b110;
        rom_memory[13435] = 3'b110;
        rom_memory[13436] = 3'b110;
        rom_memory[13437] = 3'b110;
        rom_memory[13438] = 3'b110;
        rom_memory[13439] = 3'b110;
        rom_memory[13440] = 3'b110;
        rom_memory[13441] = 3'b110;
        rom_memory[13442] = 3'b110;
        rom_memory[13443] = 3'b110;
        rom_memory[13444] = 3'b110;
        rom_memory[13445] = 3'b110;
        rom_memory[13446] = 3'b110;
        rom_memory[13447] = 3'b110;
        rom_memory[13448] = 3'b110;
        rom_memory[13449] = 3'b110;
        rom_memory[13450] = 3'b110;
        rom_memory[13451] = 3'b110;
        rom_memory[13452] = 3'b110;
        rom_memory[13453] = 3'b110;
        rom_memory[13454] = 3'b110;
        rom_memory[13455] = 3'b110;
        rom_memory[13456] = 3'b110;
        rom_memory[13457] = 3'b110;
        rom_memory[13458] = 3'b110;
        rom_memory[13459] = 3'b110;
        rom_memory[13460] = 3'b110;
        rom_memory[13461] = 3'b110;
        rom_memory[13462] = 3'b110;
        rom_memory[13463] = 3'b110;
        rom_memory[13464] = 3'b110;
        rom_memory[13465] = 3'b110;
        rom_memory[13466] = 3'b110;
        rom_memory[13467] = 3'b110;
        rom_memory[13468] = 3'b110;
        rom_memory[13469] = 3'b110;
        rom_memory[13470] = 3'b110;
        rom_memory[13471] = 3'b110;
        rom_memory[13472] = 3'b110;
        rom_memory[13473] = 3'b110;
        rom_memory[13474] = 3'b110;
        rom_memory[13475] = 3'b110;
        rom_memory[13476] = 3'b110;
        rom_memory[13477] = 3'b110;
        rom_memory[13478] = 3'b111;
        rom_memory[13479] = 3'b111;
        rom_memory[13480] = 3'b111;
        rom_memory[13481] = 3'b111;
        rom_memory[13482] = 3'b111;
        rom_memory[13483] = 3'b111;
        rom_memory[13484] = 3'b111;
        rom_memory[13485] = 3'b111;
        rom_memory[13486] = 3'b111;
        rom_memory[13487] = 3'b111;
        rom_memory[13488] = 3'b001;
        rom_memory[13489] = 3'b000;
        rom_memory[13490] = 3'b000;
        rom_memory[13491] = 3'b000;
        rom_memory[13492] = 3'b000;
        rom_memory[13493] = 3'b000;
        rom_memory[13494] = 3'b000;
        rom_memory[13495] = 3'b000;
        rom_memory[13496] = 3'b000;
        rom_memory[13497] = 3'b000;
        rom_memory[13498] = 3'b000;
        rom_memory[13499] = 3'b000;
        rom_memory[13500] = 3'b000;
        rom_memory[13501] = 3'b000;
        rom_memory[13502] = 3'b000;
        rom_memory[13503] = 3'b000;
        rom_memory[13504] = 3'b000;
        rom_memory[13505] = 3'b000;
        rom_memory[13506] = 3'b000;
        rom_memory[13507] = 3'b000;
        rom_memory[13508] = 3'b000;
        rom_memory[13509] = 3'b000;
        rom_memory[13510] = 3'b000;
        rom_memory[13511] = 3'b000;
        rom_memory[13512] = 3'b000;
        rom_memory[13513] = 3'b000;
        rom_memory[13514] = 3'b000;
        rom_memory[13515] = 3'b000;
        rom_memory[13516] = 3'b000;
        rom_memory[13517] = 3'b000;
        rom_memory[13518] = 3'b000;
        rom_memory[13519] = 3'b000;
        rom_memory[13520] = 3'b000;
        rom_memory[13521] = 3'b001;
        rom_memory[13522] = 3'b011;
        rom_memory[13523] = 3'b011;
        rom_memory[13524] = 3'b011;
        rom_memory[13525] = 3'b011;
        rom_memory[13526] = 3'b011;
        rom_memory[13527] = 3'b011;
        rom_memory[13528] = 3'b011;
        rom_memory[13529] = 3'b011;
        rom_memory[13530] = 3'b011;
        rom_memory[13531] = 3'b011;
        rom_memory[13532] = 3'b111;
        rom_memory[13533] = 3'b111;
        rom_memory[13534] = 3'b110;
        rom_memory[13535] = 3'b110;
        rom_memory[13536] = 3'b110;
        rom_memory[13537] = 3'b111;
        rom_memory[13538] = 3'b111;
        rom_memory[13539] = 3'b111;
        rom_memory[13540] = 3'b111;
        rom_memory[13541] = 3'b111;
        rom_memory[13542] = 3'b011;
        rom_memory[13543] = 3'b011;
        rom_memory[13544] = 3'b111;
        rom_memory[13545] = 3'b110;
        rom_memory[13546] = 3'b110;
        rom_memory[13547] = 3'b110;
        rom_memory[13548] = 3'b110;
        rom_memory[13549] = 3'b110;
        rom_memory[13550] = 3'b110;
        rom_memory[13551] = 3'b110;
        rom_memory[13552] = 3'b110;
        rom_memory[13553] = 3'b110;
        rom_memory[13554] = 3'b110;
        rom_memory[13555] = 3'b110;
        rom_memory[13556] = 3'b110;
        rom_memory[13557] = 3'b110;
        rom_memory[13558] = 3'b110;
        rom_memory[13559] = 3'b110;
        rom_memory[13560] = 3'b110;
        rom_memory[13561] = 3'b110;
        rom_memory[13562] = 3'b110;
        rom_memory[13563] = 3'b110;
        rom_memory[13564] = 3'b110;
        rom_memory[13565] = 3'b110;
        rom_memory[13566] = 3'b111;
        rom_memory[13567] = 3'b111;
        rom_memory[13568] = 3'b111;
        rom_memory[13569] = 3'b110;
        rom_memory[13570] = 3'b110;
        rom_memory[13571] = 3'b111;
        rom_memory[13572] = 3'b111;
        rom_memory[13573] = 3'b111;
        rom_memory[13574] = 3'b111;
        rom_memory[13575] = 3'b110;
        rom_memory[13576] = 3'b111;
        rom_memory[13577] = 3'b111;
        rom_memory[13578] = 3'b111;
        rom_memory[13579] = 3'b111;
        rom_memory[13580] = 3'b111;
        rom_memory[13581] = 3'b110;
        rom_memory[13582] = 3'b111;
        rom_memory[13583] = 3'b111;
        rom_memory[13584] = 3'b111;
        rom_memory[13585] = 3'b111;
        rom_memory[13586] = 3'b111;
        rom_memory[13587] = 3'b111;
        rom_memory[13588] = 3'b110;
        rom_memory[13589] = 3'b110;
        rom_memory[13590] = 3'b111;
        rom_memory[13591] = 3'b111;
        rom_memory[13592] = 3'b111;
        rom_memory[13593] = 3'b111;
        rom_memory[13594] = 3'b110;
        rom_memory[13595] = 3'b110;
        rom_memory[13596] = 3'b110;
        rom_memory[13597] = 3'b110;
        rom_memory[13598] = 3'b110;
        rom_memory[13599] = 3'b110;
        rom_memory[13600] = 3'b110;
        rom_memory[13601] = 3'b110;
        rom_memory[13602] = 3'b110;
        rom_memory[13603] = 3'b110;
        rom_memory[13604] = 3'b110;
        rom_memory[13605] = 3'b110;
        rom_memory[13606] = 3'b110;
        rom_memory[13607] = 3'b110;
        rom_memory[13608] = 3'b110;
        rom_memory[13609] = 3'b110;
        rom_memory[13610] = 3'b110;
        rom_memory[13611] = 3'b110;
        rom_memory[13612] = 3'b110;
        rom_memory[13613] = 3'b110;
        rom_memory[13614] = 3'b110;
        rom_memory[13615] = 3'b110;
        rom_memory[13616] = 3'b110;
        rom_memory[13617] = 3'b110;
        rom_memory[13618] = 3'b110;
        rom_memory[13619] = 3'b110;
        rom_memory[13620] = 3'b110;
        rom_memory[13621] = 3'b110;
        rom_memory[13622] = 3'b110;
        rom_memory[13623] = 3'b110;
        rom_memory[13624] = 3'b110;
        rom_memory[13625] = 3'b110;
        rom_memory[13626] = 3'b110;
        rom_memory[13627] = 3'b110;
        rom_memory[13628] = 3'b110;
        rom_memory[13629] = 3'b110;
        rom_memory[13630] = 3'b110;
        rom_memory[13631] = 3'b110;
        rom_memory[13632] = 3'b110;
        rom_memory[13633] = 3'b110;
        rom_memory[13634] = 3'b110;
        rom_memory[13635] = 3'b110;
        rom_memory[13636] = 3'b110;
        rom_memory[13637] = 3'b110;
        rom_memory[13638] = 3'b110;
        rom_memory[13639] = 3'b110;
        rom_memory[13640] = 3'b110;
        rom_memory[13641] = 3'b110;
        rom_memory[13642] = 3'b110;
        rom_memory[13643] = 3'b110;
        rom_memory[13644] = 3'b110;
        rom_memory[13645] = 3'b110;
        rom_memory[13646] = 3'b110;
        rom_memory[13647] = 3'b110;
        rom_memory[13648] = 3'b110;
        rom_memory[13649] = 3'b110;
        rom_memory[13650] = 3'b110;
        rom_memory[13651] = 3'b110;
        rom_memory[13652] = 3'b110;
        rom_memory[13653] = 3'b110;
        rom_memory[13654] = 3'b110;
        rom_memory[13655] = 3'b110;
        rom_memory[13656] = 3'b110;
        rom_memory[13657] = 3'b110;
        rom_memory[13658] = 3'b110;
        rom_memory[13659] = 3'b110;
        rom_memory[13660] = 3'b110;
        rom_memory[13661] = 3'b110;
        rom_memory[13662] = 3'b110;
        rom_memory[13663] = 3'b110;
        rom_memory[13664] = 3'b110;
        rom_memory[13665] = 3'b110;
        rom_memory[13666] = 3'b110;
        rom_memory[13667] = 3'b110;
        rom_memory[13668] = 3'b110;
        rom_memory[13669] = 3'b110;
        rom_memory[13670] = 3'b110;
        rom_memory[13671] = 3'b110;
        rom_memory[13672] = 3'b110;
        rom_memory[13673] = 3'b110;
        rom_memory[13674] = 3'b110;
        rom_memory[13675] = 3'b110;
        rom_memory[13676] = 3'b110;
        rom_memory[13677] = 3'b110;
        rom_memory[13678] = 3'b110;
        rom_memory[13679] = 3'b110;
        rom_memory[13680] = 3'b110;
        rom_memory[13681] = 3'b110;
        rom_memory[13682] = 3'b110;
        rom_memory[13683] = 3'b110;
        rom_memory[13684] = 3'b110;
        rom_memory[13685] = 3'b110;
        rom_memory[13686] = 3'b110;
        rom_memory[13687] = 3'b110;
        rom_memory[13688] = 3'b110;
        rom_memory[13689] = 3'b110;
        rom_memory[13690] = 3'b110;
        rom_memory[13691] = 3'b110;
        rom_memory[13692] = 3'b110;
        rom_memory[13693] = 3'b110;
        rom_memory[13694] = 3'b110;
        rom_memory[13695] = 3'b110;
        rom_memory[13696] = 3'b110;
        rom_memory[13697] = 3'b110;
        rom_memory[13698] = 3'b110;
        rom_memory[13699] = 3'b110;
        rom_memory[13700] = 3'b110;
        rom_memory[13701] = 3'b110;
        rom_memory[13702] = 3'b110;
        rom_memory[13703] = 3'b110;
        rom_memory[13704] = 3'b110;
        rom_memory[13705] = 3'b110;
        rom_memory[13706] = 3'b110;
        rom_memory[13707] = 3'b110;
        rom_memory[13708] = 3'b110;
        rom_memory[13709] = 3'b110;
        rom_memory[13710] = 3'b110;
        rom_memory[13711] = 3'b110;
        rom_memory[13712] = 3'b110;
        rom_memory[13713] = 3'b110;
        rom_memory[13714] = 3'b110;
        rom_memory[13715] = 3'b110;
        rom_memory[13716] = 3'b110;
        rom_memory[13717] = 3'b110;
        rom_memory[13718] = 3'b111;
        rom_memory[13719] = 3'b111;
        rom_memory[13720] = 3'b111;
        rom_memory[13721] = 3'b111;
        rom_memory[13722] = 3'b111;
        rom_memory[13723] = 3'b111;
        rom_memory[13724] = 3'b111;
        rom_memory[13725] = 3'b111;
        rom_memory[13726] = 3'b111;
        rom_memory[13727] = 3'b111;
        rom_memory[13728] = 3'b000;
        rom_memory[13729] = 3'b000;
        rom_memory[13730] = 3'b000;
        rom_memory[13731] = 3'b000;
        rom_memory[13732] = 3'b000;
        rom_memory[13733] = 3'b000;
        rom_memory[13734] = 3'b000;
        rom_memory[13735] = 3'b000;
        rom_memory[13736] = 3'b000;
        rom_memory[13737] = 3'b000;
        rom_memory[13738] = 3'b000;
        rom_memory[13739] = 3'b000;
        rom_memory[13740] = 3'b000;
        rom_memory[13741] = 3'b000;
        rom_memory[13742] = 3'b000;
        rom_memory[13743] = 3'b000;
        rom_memory[13744] = 3'b000;
        rom_memory[13745] = 3'b000;
        rom_memory[13746] = 3'b000;
        rom_memory[13747] = 3'b000;
        rom_memory[13748] = 3'b000;
        rom_memory[13749] = 3'b000;
        rom_memory[13750] = 3'b000;
        rom_memory[13751] = 3'b000;
        rom_memory[13752] = 3'b000;
        rom_memory[13753] = 3'b000;
        rom_memory[13754] = 3'b000;
        rom_memory[13755] = 3'b000;
        rom_memory[13756] = 3'b000;
        rom_memory[13757] = 3'b000;
        rom_memory[13758] = 3'b000;
        rom_memory[13759] = 3'b000;
        rom_memory[13760] = 3'b000;
        rom_memory[13761] = 3'b000;
        rom_memory[13762] = 3'b011;
        rom_memory[13763] = 3'b011;
        rom_memory[13764] = 3'b011;
        rom_memory[13765] = 3'b011;
        rom_memory[13766] = 3'b011;
        rom_memory[13767] = 3'b011;
        rom_memory[13768] = 3'b011;
        rom_memory[13769] = 3'b011;
        rom_memory[13770] = 3'b011;
        rom_memory[13771] = 3'b011;
        rom_memory[13772] = 3'b111;
        rom_memory[13773] = 3'b111;
        rom_memory[13774] = 3'b110;
        rom_memory[13775] = 3'b110;
        rom_memory[13776] = 3'b110;
        rom_memory[13777] = 3'b110;
        rom_memory[13778] = 3'b111;
        rom_memory[13779] = 3'b111;
        rom_memory[13780] = 3'b111;
        rom_memory[13781] = 3'b111;
        rom_memory[13782] = 3'b111;
        rom_memory[13783] = 3'b111;
        rom_memory[13784] = 3'b111;
        rom_memory[13785] = 3'b110;
        rom_memory[13786] = 3'b110;
        rom_memory[13787] = 3'b110;
        rom_memory[13788] = 3'b110;
        rom_memory[13789] = 3'b110;
        rom_memory[13790] = 3'b110;
        rom_memory[13791] = 3'b110;
        rom_memory[13792] = 3'b110;
        rom_memory[13793] = 3'b110;
        rom_memory[13794] = 3'b110;
        rom_memory[13795] = 3'b110;
        rom_memory[13796] = 3'b110;
        rom_memory[13797] = 3'b110;
        rom_memory[13798] = 3'b110;
        rom_memory[13799] = 3'b110;
        rom_memory[13800] = 3'b110;
        rom_memory[13801] = 3'b110;
        rom_memory[13802] = 3'b110;
        rom_memory[13803] = 3'b110;
        rom_memory[13804] = 3'b110;
        rom_memory[13805] = 3'b110;
        rom_memory[13806] = 3'b111;
        rom_memory[13807] = 3'b111;
        rom_memory[13808] = 3'b111;
        rom_memory[13809] = 3'b111;
        rom_memory[13810] = 3'b111;
        rom_memory[13811] = 3'b111;
        rom_memory[13812] = 3'b111;
        rom_memory[13813] = 3'b110;
        rom_memory[13814] = 3'b111;
        rom_memory[13815] = 3'b111;
        rom_memory[13816] = 3'b111;
        rom_memory[13817] = 3'b111;
        rom_memory[13818] = 3'b110;
        rom_memory[13819] = 3'b110;
        rom_memory[13820] = 3'b111;
        rom_memory[13821] = 3'b111;
        rom_memory[13822] = 3'b111;
        rom_memory[13823] = 3'b111;
        rom_memory[13824] = 3'b111;
        rom_memory[13825] = 3'b111;
        rom_memory[13826] = 3'b111;
        rom_memory[13827] = 3'b111;
        rom_memory[13828] = 3'b111;
        rom_memory[13829] = 3'b111;
        rom_memory[13830] = 3'b110;
        rom_memory[13831] = 3'b111;
        rom_memory[13832] = 3'b111;
        rom_memory[13833] = 3'b111;
        rom_memory[13834] = 3'b111;
        rom_memory[13835] = 3'b111;
        rom_memory[13836] = 3'b111;
        rom_memory[13837] = 3'b110;
        rom_memory[13838] = 3'b110;
        rom_memory[13839] = 3'b110;
        rom_memory[13840] = 3'b110;
        rom_memory[13841] = 3'b110;
        rom_memory[13842] = 3'b110;
        rom_memory[13843] = 3'b110;
        rom_memory[13844] = 3'b110;
        rom_memory[13845] = 3'b110;
        rom_memory[13846] = 3'b110;
        rom_memory[13847] = 3'b110;
        rom_memory[13848] = 3'b110;
        rom_memory[13849] = 3'b110;
        rom_memory[13850] = 3'b110;
        rom_memory[13851] = 3'b110;
        rom_memory[13852] = 3'b110;
        rom_memory[13853] = 3'b110;
        rom_memory[13854] = 3'b110;
        rom_memory[13855] = 3'b110;
        rom_memory[13856] = 3'b110;
        rom_memory[13857] = 3'b110;
        rom_memory[13858] = 3'b110;
        rom_memory[13859] = 3'b110;
        rom_memory[13860] = 3'b110;
        rom_memory[13861] = 3'b110;
        rom_memory[13862] = 3'b110;
        rom_memory[13863] = 3'b110;
        rom_memory[13864] = 3'b110;
        rom_memory[13865] = 3'b110;
        rom_memory[13866] = 3'b110;
        rom_memory[13867] = 3'b110;
        rom_memory[13868] = 3'b110;
        rom_memory[13869] = 3'b110;
        rom_memory[13870] = 3'b110;
        rom_memory[13871] = 3'b110;
        rom_memory[13872] = 3'b110;
        rom_memory[13873] = 3'b110;
        rom_memory[13874] = 3'b110;
        rom_memory[13875] = 3'b110;
        rom_memory[13876] = 3'b110;
        rom_memory[13877] = 3'b110;
        rom_memory[13878] = 3'b110;
        rom_memory[13879] = 3'b110;
        rom_memory[13880] = 3'b110;
        rom_memory[13881] = 3'b110;
        rom_memory[13882] = 3'b110;
        rom_memory[13883] = 3'b110;
        rom_memory[13884] = 3'b110;
        rom_memory[13885] = 3'b110;
        rom_memory[13886] = 3'b110;
        rom_memory[13887] = 3'b110;
        rom_memory[13888] = 3'b110;
        rom_memory[13889] = 3'b110;
        rom_memory[13890] = 3'b110;
        rom_memory[13891] = 3'b110;
        rom_memory[13892] = 3'b110;
        rom_memory[13893] = 3'b110;
        rom_memory[13894] = 3'b110;
        rom_memory[13895] = 3'b110;
        rom_memory[13896] = 3'b110;
        rom_memory[13897] = 3'b110;
        rom_memory[13898] = 3'b110;
        rom_memory[13899] = 3'b110;
        rom_memory[13900] = 3'b110;
        rom_memory[13901] = 3'b110;
        rom_memory[13902] = 3'b110;
        rom_memory[13903] = 3'b110;
        rom_memory[13904] = 3'b110;
        rom_memory[13905] = 3'b110;
        rom_memory[13906] = 3'b110;
        rom_memory[13907] = 3'b110;
        rom_memory[13908] = 3'b110;
        rom_memory[13909] = 3'b110;
        rom_memory[13910] = 3'b110;
        rom_memory[13911] = 3'b110;
        rom_memory[13912] = 3'b110;
        rom_memory[13913] = 3'b110;
        rom_memory[13914] = 3'b110;
        rom_memory[13915] = 3'b110;
        rom_memory[13916] = 3'b110;
        rom_memory[13917] = 3'b110;
        rom_memory[13918] = 3'b110;
        rom_memory[13919] = 3'b110;
        rom_memory[13920] = 3'b110;
        rom_memory[13921] = 3'b110;
        rom_memory[13922] = 3'b110;
        rom_memory[13923] = 3'b110;
        rom_memory[13924] = 3'b110;
        rom_memory[13925] = 3'b110;
        rom_memory[13926] = 3'b110;
        rom_memory[13927] = 3'b110;
        rom_memory[13928] = 3'b110;
        rom_memory[13929] = 3'b110;
        rom_memory[13930] = 3'b110;
        rom_memory[13931] = 3'b110;
        rom_memory[13932] = 3'b110;
        rom_memory[13933] = 3'b110;
        rom_memory[13934] = 3'b110;
        rom_memory[13935] = 3'b110;
        rom_memory[13936] = 3'b110;
        rom_memory[13937] = 3'b110;
        rom_memory[13938] = 3'b110;
        rom_memory[13939] = 3'b110;
        rom_memory[13940] = 3'b110;
        rom_memory[13941] = 3'b110;
        rom_memory[13942] = 3'b110;
        rom_memory[13943] = 3'b110;
        rom_memory[13944] = 3'b110;
        rom_memory[13945] = 3'b110;
        rom_memory[13946] = 3'b110;
        rom_memory[13947] = 3'b110;
        rom_memory[13948] = 3'b110;
        rom_memory[13949] = 3'b110;
        rom_memory[13950] = 3'b110;
        rom_memory[13951] = 3'b110;
        rom_memory[13952] = 3'b110;
        rom_memory[13953] = 3'b110;
        rom_memory[13954] = 3'b110;
        rom_memory[13955] = 3'b110;
        rom_memory[13956] = 3'b110;
        rom_memory[13957] = 3'b111;
        rom_memory[13958] = 3'b111;
        rom_memory[13959] = 3'b111;
        rom_memory[13960] = 3'b111;
        rom_memory[13961] = 3'b111;
        rom_memory[13962] = 3'b111;
        rom_memory[13963] = 3'b111;
        rom_memory[13964] = 3'b111;
        rom_memory[13965] = 3'b111;
        rom_memory[13966] = 3'b111;
        rom_memory[13967] = 3'b111;
        rom_memory[13968] = 3'b000;
        rom_memory[13969] = 3'b000;
        rom_memory[13970] = 3'b000;
        rom_memory[13971] = 3'b000;
        rom_memory[13972] = 3'b000;
        rom_memory[13973] = 3'b000;
        rom_memory[13974] = 3'b000;
        rom_memory[13975] = 3'b000;
        rom_memory[13976] = 3'b000;
        rom_memory[13977] = 3'b000;
        rom_memory[13978] = 3'b000;
        rom_memory[13979] = 3'b000;
        rom_memory[13980] = 3'b000;
        rom_memory[13981] = 3'b000;
        rom_memory[13982] = 3'b000;
        rom_memory[13983] = 3'b000;
        rom_memory[13984] = 3'b000;
        rom_memory[13985] = 3'b000;
        rom_memory[13986] = 3'b000;
        rom_memory[13987] = 3'b000;
        rom_memory[13988] = 3'b000;
        rom_memory[13989] = 3'b000;
        rom_memory[13990] = 3'b000;
        rom_memory[13991] = 3'b000;
        rom_memory[13992] = 3'b000;
        rom_memory[13993] = 3'b000;
        rom_memory[13994] = 3'b000;
        rom_memory[13995] = 3'b000;
        rom_memory[13996] = 3'b000;
        rom_memory[13997] = 3'b000;
        rom_memory[13998] = 3'b000;
        rom_memory[13999] = 3'b000;
        rom_memory[14000] = 3'b111;
        rom_memory[14001] = 3'b000;
        rom_memory[14002] = 3'b000;
        rom_memory[14003] = 3'b000;
        rom_memory[14004] = 3'b011;
        rom_memory[14005] = 3'b011;
        rom_memory[14006] = 3'b011;
        rom_memory[14007] = 3'b011;
        rom_memory[14008] = 3'b011;
        rom_memory[14009] = 3'b111;
        rom_memory[14010] = 3'b011;
        rom_memory[14011] = 3'b011;
        rom_memory[14012] = 3'b011;
        rom_memory[14013] = 3'b110;
        rom_memory[14014] = 3'b110;
        rom_memory[14015] = 3'b110;
        rom_memory[14016] = 3'b110;
        rom_memory[14017] = 3'b110;
        rom_memory[14018] = 3'b110;
        rom_memory[14019] = 3'b111;
        rom_memory[14020] = 3'b111;
        rom_memory[14021] = 3'b111;
        rom_memory[14022] = 3'b111;
        rom_memory[14023] = 3'b111;
        rom_memory[14024] = 3'b110;
        rom_memory[14025] = 3'b110;
        rom_memory[14026] = 3'b110;
        rom_memory[14027] = 3'b110;
        rom_memory[14028] = 3'b110;
        rom_memory[14029] = 3'b110;
        rom_memory[14030] = 3'b110;
        rom_memory[14031] = 3'b110;
        rom_memory[14032] = 3'b110;
        rom_memory[14033] = 3'b110;
        rom_memory[14034] = 3'b110;
        rom_memory[14035] = 3'b110;
        rom_memory[14036] = 3'b110;
        rom_memory[14037] = 3'b110;
        rom_memory[14038] = 3'b110;
        rom_memory[14039] = 3'b110;
        rom_memory[14040] = 3'b110;
        rom_memory[14041] = 3'b110;
        rom_memory[14042] = 3'b110;
        rom_memory[14043] = 3'b110;
        rom_memory[14044] = 3'b110;
        rom_memory[14045] = 3'b110;
        rom_memory[14046] = 3'b111;
        rom_memory[14047] = 3'b111;
        rom_memory[14048] = 3'b111;
        rom_memory[14049] = 3'b111;
        rom_memory[14050] = 3'b111;
        rom_memory[14051] = 3'b111;
        rom_memory[14052] = 3'b111;
        rom_memory[14053] = 3'b111;
        rom_memory[14054] = 3'b111;
        rom_memory[14055] = 3'b111;
        rom_memory[14056] = 3'b111;
        rom_memory[14057] = 3'b111;
        rom_memory[14058] = 3'b111;
        rom_memory[14059] = 3'b111;
        rom_memory[14060] = 3'b111;
        rom_memory[14061] = 3'b111;
        rom_memory[14062] = 3'b111;
        rom_memory[14063] = 3'b111;
        rom_memory[14064] = 3'b111;
        rom_memory[14065] = 3'b111;
        rom_memory[14066] = 3'b111;
        rom_memory[14067] = 3'b111;
        rom_memory[14068] = 3'b111;
        rom_memory[14069] = 3'b110;
        rom_memory[14070] = 3'b111;
        rom_memory[14071] = 3'b111;
        rom_memory[14072] = 3'b111;
        rom_memory[14073] = 3'b111;
        rom_memory[14074] = 3'b111;
        rom_memory[14075] = 3'b111;
        rom_memory[14076] = 3'b111;
        rom_memory[14077] = 3'b110;
        rom_memory[14078] = 3'b110;
        rom_memory[14079] = 3'b110;
        rom_memory[14080] = 3'b110;
        rom_memory[14081] = 3'b110;
        rom_memory[14082] = 3'b110;
        rom_memory[14083] = 3'b110;
        rom_memory[14084] = 3'b110;
        rom_memory[14085] = 3'b110;
        rom_memory[14086] = 3'b110;
        rom_memory[14087] = 3'b110;
        rom_memory[14088] = 3'b110;
        rom_memory[14089] = 3'b110;
        rom_memory[14090] = 3'b110;
        rom_memory[14091] = 3'b110;
        rom_memory[14092] = 3'b110;
        rom_memory[14093] = 3'b110;
        rom_memory[14094] = 3'b110;
        rom_memory[14095] = 3'b110;
        rom_memory[14096] = 3'b110;
        rom_memory[14097] = 3'b110;
        rom_memory[14098] = 3'b110;
        rom_memory[14099] = 3'b110;
        rom_memory[14100] = 3'b110;
        rom_memory[14101] = 3'b110;
        rom_memory[14102] = 3'b110;
        rom_memory[14103] = 3'b110;
        rom_memory[14104] = 3'b110;
        rom_memory[14105] = 3'b110;
        rom_memory[14106] = 3'b110;
        rom_memory[14107] = 3'b110;
        rom_memory[14108] = 3'b110;
        rom_memory[14109] = 3'b110;
        rom_memory[14110] = 3'b110;
        rom_memory[14111] = 3'b110;
        rom_memory[14112] = 3'b110;
        rom_memory[14113] = 3'b110;
        rom_memory[14114] = 3'b110;
        rom_memory[14115] = 3'b110;
        rom_memory[14116] = 3'b110;
        rom_memory[14117] = 3'b110;
        rom_memory[14118] = 3'b110;
        rom_memory[14119] = 3'b110;
        rom_memory[14120] = 3'b110;
        rom_memory[14121] = 3'b110;
        rom_memory[14122] = 3'b110;
        rom_memory[14123] = 3'b110;
        rom_memory[14124] = 3'b110;
        rom_memory[14125] = 3'b110;
        rom_memory[14126] = 3'b110;
        rom_memory[14127] = 3'b110;
        rom_memory[14128] = 3'b110;
        rom_memory[14129] = 3'b110;
        rom_memory[14130] = 3'b110;
        rom_memory[14131] = 3'b110;
        rom_memory[14132] = 3'b110;
        rom_memory[14133] = 3'b110;
        rom_memory[14134] = 3'b110;
        rom_memory[14135] = 3'b110;
        rom_memory[14136] = 3'b110;
        rom_memory[14137] = 3'b110;
        rom_memory[14138] = 3'b110;
        rom_memory[14139] = 3'b110;
        rom_memory[14140] = 3'b110;
        rom_memory[14141] = 3'b110;
        rom_memory[14142] = 3'b110;
        rom_memory[14143] = 3'b110;
        rom_memory[14144] = 3'b110;
        rom_memory[14145] = 3'b110;
        rom_memory[14146] = 3'b110;
        rom_memory[14147] = 3'b110;
        rom_memory[14148] = 3'b110;
        rom_memory[14149] = 3'b110;
        rom_memory[14150] = 3'b110;
        rom_memory[14151] = 3'b110;
        rom_memory[14152] = 3'b110;
        rom_memory[14153] = 3'b110;
        rom_memory[14154] = 3'b110;
        rom_memory[14155] = 3'b110;
        rom_memory[14156] = 3'b110;
        rom_memory[14157] = 3'b110;
        rom_memory[14158] = 3'b110;
        rom_memory[14159] = 3'b110;
        rom_memory[14160] = 3'b110;
        rom_memory[14161] = 3'b110;
        rom_memory[14162] = 3'b110;
        rom_memory[14163] = 3'b110;
        rom_memory[14164] = 3'b110;
        rom_memory[14165] = 3'b110;
        rom_memory[14166] = 3'b110;
        rom_memory[14167] = 3'b110;
        rom_memory[14168] = 3'b110;
        rom_memory[14169] = 3'b110;
        rom_memory[14170] = 3'b110;
        rom_memory[14171] = 3'b110;
        rom_memory[14172] = 3'b110;
        rom_memory[14173] = 3'b110;
        rom_memory[14174] = 3'b110;
        rom_memory[14175] = 3'b110;
        rom_memory[14176] = 3'b110;
        rom_memory[14177] = 3'b110;
        rom_memory[14178] = 3'b110;
        rom_memory[14179] = 3'b110;
        rom_memory[14180] = 3'b110;
        rom_memory[14181] = 3'b110;
        rom_memory[14182] = 3'b110;
        rom_memory[14183] = 3'b110;
        rom_memory[14184] = 3'b110;
        rom_memory[14185] = 3'b110;
        rom_memory[14186] = 3'b110;
        rom_memory[14187] = 3'b110;
        rom_memory[14188] = 3'b110;
        rom_memory[14189] = 3'b110;
        rom_memory[14190] = 3'b110;
        rom_memory[14191] = 3'b110;
        rom_memory[14192] = 3'b110;
        rom_memory[14193] = 3'b110;
        rom_memory[14194] = 3'b110;
        rom_memory[14195] = 3'b110;
        rom_memory[14196] = 3'b110;
        rom_memory[14197] = 3'b110;
        rom_memory[14198] = 3'b111;
        rom_memory[14199] = 3'b111;
        rom_memory[14200] = 3'b111;
        rom_memory[14201] = 3'b111;
        rom_memory[14202] = 3'b111;
        rom_memory[14203] = 3'b111;
        rom_memory[14204] = 3'b111;
        rom_memory[14205] = 3'b111;
        rom_memory[14206] = 3'b111;
        rom_memory[14207] = 3'b001;
        rom_memory[14208] = 3'b000;
        rom_memory[14209] = 3'b000;
        rom_memory[14210] = 3'b000;
        rom_memory[14211] = 3'b000;
        rom_memory[14212] = 3'b000;
        rom_memory[14213] = 3'b000;
        rom_memory[14214] = 3'b000;
        rom_memory[14215] = 3'b000;
        rom_memory[14216] = 3'b000;
        rom_memory[14217] = 3'b000;
        rom_memory[14218] = 3'b000;
        rom_memory[14219] = 3'b000;
        rom_memory[14220] = 3'b000;
        rom_memory[14221] = 3'b000;
        rom_memory[14222] = 3'b000;
        rom_memory[14223] = 3'b000;
        rom_memory[14224] = 3'b000;
        rom_memory[14225] = 3'b000;
        rom_memory[14226] = 3'b000;
        rom_memory[14227] = 3'b000;
        rom_memory[14228] = 3'b000;
        rom_memory[14229] = 3'b000;
        rom_memory[14230] = 3'b000;
        rom_memory[14231] = 3'b000;
        rom_memory[14232] = 3'b000;
        rom_memory[14233] = 3'b000;
        rom_memory[14234] = 3'b000;
        rom_memory[14235] = 3'b000;
        rom_memory[14236] = 3'b000;
        rom_memory[14237] = 3'b000;
        rom_memory[14238] = 3'b000;
        rom_memory[14239] = 3'b100;
        rom_memory[14240] = 3'b111;
        rom_memory[14241] = 3'b110;
        rom_memory[14242] = 3'b000;
        rom_memory[14243] = 3'b000;
        rom_memory[14244] = 3'b001;
        rom_memory[14245] = 3'b011;
        rom_memory[14246] = 3'b011;
        rom_memory[14247] = 3'b011;
        rom_memory[14248] = 3'b011;
        rom_memory[14249] = 3'b011;
        rom_memory[14250] = 3'b011;
        rom_memory[14251] = 3'b011;
        rom_memory[14252] = 3'b111;
        rom_memory[14253] = 3'b110;
        rom_memory[14254] = 3'b110;
        rom_memory[14255] = 3'b110;
        rom_memory[14256] = 3'b110;
        rom_memory[14257] = 3'b110;
        rom_memory[14258] = 3'b110;
        rom_memory[14259] = 3'b111;
        rom_memory[14260] = 3'b111;
        rom_memory[14261] = 3'b110;
        rom_memory[14262] = 3'b110;
        rom_memory[14263] = 3'b111;
        rom_memory[14264] = 3'b111;
        rom_memory[14265] = 3'b110;
        rom_memory[14266] = 3'b110;
        rom_memory[14267] = 3'b110;
        rom_memory[14268] = 3'b110;
        rom_memory[14269] = 3'b110;
        rom_memory[14270] = 3'b110;
        rom_memory[14271] = 3'b110;
        rom_memory[14272] = 3'b110;
        rom_memory[14273] = 3'b110;
        rom_memory[14274] = 3'b110;
        rom_memory[14275] = 3'b110;
        rom_memory[14276] = 3'b110;
        rom_memory[14277] = 3'b110;
        rom_memory[14278] = 3'b110;
        rom_memory[14279] = 3'b110;
        rom_memory[14280] = 3'b110;
        rom_memory[14281] = 3'b110;
        rom_memory[14282] = 3'b110;
        rom_memory[14283] = 3'b110;
        rom_memory[14284] = 3'b110;
        rom_memory[14285] = 3'b110;
        rom_memory[14286] = 3'b110;
        rom_memory[14287] = 3'b110;
        rom_memory[14288] = 3'b110;
        rom_memory[14289] = 3'b110;
        rom_memory[14290] = 3'b111;
        rom_memory[14291] = 3'b111;
        rom_memory[14292] = 3'b111;
        rom_memory[14293] = 3'b111;
        rom_memory[14294] = 3'b111;
        rom_memory[14295] = 3'b111;
        rom_memory[14296] = 3'b111;
        rom_memory[14297] = 3'b111;
        rom_memory[14298] = 3'b111;
        rom_memory[14299] = 3'b111;
        rom_memory[14300] = 3'b111;
        rom_memory[14301] = 3'b111;
        rom_memory[14302] = 3'b111;
        rom_memory[14303] = 3'b111;
        rom_memory[14304] = 3'b111;
        rom_memory[14305] = 3'b111;
        rom_memory[14306] = 3'b111;
        rom_memory[14307] = 3'b111;
        rom_memory[14308] = 3'b111;
        rom_memory[14309] = 3'b111;
        rom_memory[14310] = 3'b111;
        rom_memory[14311] = 3'b111;
        rom_memory[14312] = 3'b111;
        rom_memory[14313] = 3'b111;
        rom_memory[14314] = 3'b111;
        rom_memory[14315] = 3'b110;
        rom_memory[14316] = 3'b111;
        rom_memory[14317] = 3'b111;
        rom_memory[14318] = 3'b110;
        rom_memory[14319] = 3'b110;
        rom_memory[14320] = 3'b110;
        rom_memory[14321] = 3'b110;
        rom_memory[14322] = 3'b110;
        rom_memory[14323] = 3'b110;
        rom_memory[14324] = 3'b110;
        rom_memory[14325] = 3'b110;
        rom_memory[14326] = 3'b110;
        rom_memory[14327] = 3'b110;
        rom_memory[14328] = 3'b110;
        rom_memory[14329] = 3'b110;
        rom_memory[14330] = 3'b110;
        rom_memory[14331] = 3'b110;
        rom_memory[14332] = 3'b110;
        rom_memory[14333] = 3'b110;
        rom_memory[14334] = 3'b110;
        rom_memory[14335] = 3'b110;
        rom_memory[14336] = 3'b110;
        rom_memory[14337] = 3'b110;
        rom_memory[14338] = 3'b110;
        rom_memory[14339] = 3'b110;
        rom_memory[14340] = 3'b110;
        rom_memory[14341] = 3'b110;
        rom_memory[14342] = 3'b110;
        rom_memory[14343] = 3'b110;
        rom_memory[14344] = 3'b110;
        rom_memory[14345] = 3'b110;
        rom_memory[14346] = 3'b110;
        rom_memory[14347] = 3'b110;
        rom_memory[14348] = 3'b110;
        rom_memory[14349] = 3'b110;
        rom_memory[14350] = 3'b110;
        rom_memory[14351] = 3'b110;
        rom_memory[14352] = 3'b110;
        rom_memory[14353] = 3'b110;
        rom_memory[14354] = 3'b110;
        rom_memory[14355] = 3'b110;
        rom_memory[14356] = 3'b110;
        rom_memory[14357] = 3'b110;
        rom_memory[14358] = 3'b110;
        rom_memory[14359] = 3'b110;
        rom_memory[14360] = 3'b110;
        rom_memory[14361] = 3'b110;
        rom_memory[14362] = 3'b110;
        rom_memory[14363] = 3'b110;
        rom_memory[14364] = 3'b110;
        rom_memory[14365] = 3'b110;
        rom_memory[14366] = 3'b110;
        rom_memory[14367] = 3'b110;
        rom_memory[14368] = 3'b110;
        rom_memory[14369] = 3'b110;
        rom_memory[14370] = 3'b110;
        rom_memory[14371] = 3'b110;
        rom_memory[14372] = 3'b110;
        rom_memory[14373] = 3'b110;
        rom_memory[14374] = 3'b110;
        rom_memory[14375] = 3'b110;
        rom_memory[14376] = 3'b110;
        rom_memory[14377] = 3'b110;
        rom_memory[14378] = 3'b110;
        rom_memory[14379] = 3'b110;
        rom_memory[14380] = 3'b110;
        rom_memory[14381] = 3'b110;
        rom_memory[14382] = 3'b110;
        rom_memory[14383] = 3'b110;
        rom_memory[14384] = 3'b110;
        rom_memory[14385] = 3'b110;
        rom_memory[14386] = 3'b110;
        rom_memory[14387] = 3'b110;
        rom_memory[14388] = 3'b110;
        rom_memory[14389] = 3'b110;
        rom_memory[14390] = 3'b110;
        rom_memory[14391] = 3'b110;
        rom_memory[14392] = 3'b110;
        rom_memory[14393] = 3'b110;
        rom_memory[14394] = 3'b110;
        rom_memory[14395] = 3'b110;
        rom_memory[14396] = 3'b110;
        rom_memory[14397] = 3'b110;
        rom_memory[14398] = 3'b110;
        rom_memory[14399] = 3'b110;
        rom_memory[14400] = 3'b110;
        rom_memory[14401] = 3'b110;
        rom_memory[14402] = 3'b110;
        rom_memory[14403] = 3'b110;
        rom_memory[14404] = 3'b110;
        rom_memory[14405] = 3'b110;
        rom_memory[14406] = 3'b110;
        rom_memory[14407] = 3'b110;
        rom_memory[14408] = 3'b110;
        rom_memory[14409] = 3'b110;
        rom_memory[14410] = 3'b110;
        rom_memory[14411] = 3'b110;
        rom_memory[14412] = 3'b110;
        rom_memory[14413] = 3'b110;
        rom_memory[14414] = 3'b110;
        rom_memory[14415] = 3'b110;
        rom_memory[14416] = 3'b110;
        rom_memory[14417] = 3'b110;
        rom_memory[14418] = 3'b110;
        rom_memory[14419] = 3'b110;
        rom_memory[14420] = 3'b110;
        rom_memory[14421] = 3'b110;
        rom_memory[14422] = 3'b110;
        rom_memory[14423] = 3'b110;
        rom_memory[14424] = 3'b110;
        rom_memory[14425] = 3'b110;
        rom_memory[14426] = 3'b110;
        rom_memory[14427] = 3'b110;
        rom_memory[14428] = 3'b110;
        rom_memory[14429] = 3'b110;
        rom_memory[14430] = 3'b110;
        rom_memory[14431] = 3'b110;
        rom_memory[14432] = 3'b110;
        rom_memory[14433] = 3'b110;
        rom_memory[14434] = 3'b110;
        rom_memory[14435] = 3'b110;
        rom_memory[14436] = 3'b110;
        rom_memory[14437] = 3'b110;
        rom_memory[14438] = 3'b111;
        rom_memory[14439] = 3'b111;
        rom_memory[14440] = 3'b111;
        rom_memory[14441] = 3'b111;
        rom_memory[14442] = 3'b111;
        rom_memory[14443] = 3'b111;
        rom_memory[14444] = 3'b111;
        rom_memory[14445] = 3'b111;
        rom_memory[14446] = 3'b111;
        rom_memory[14447] = 3'b001;
        rom_memory[14448] = 3'b000;
        rom_memory[14449] = 3'b000;
        rom_memory[14450] = 3'b000;
        rom_memory[14451] = 3'b000;
        rom_memory[14452] = 3'b000;
        rom_memory[14453] = 3'b000;
        rom_memory[14454] = 3'b000;
        rom_memory[14455] = 3'b000;
        rom_memory[14456] = 3'b000;
        rom_memory[14457] = 3'b000;
        rom_memory[14458] = 3'b000;
        rom_memory[14459] = 3'b000;
        rom_memory[14460] = 3'b000;
        rom_memory[14461] = 3'b000;
        rom_memory[14462] = 3'b000;
        rom_memory[14463] = 3'b000;
        rom_memory[14464] = 3'b000;
        rom_memory[14465] = 3'b000;
        rom_memory[14466] = 3'b000;
        rom_memory[14467] = 3'b000;
        rom_memory[14468] = 3'b000;
        rom_memory[14469] = 3'b000;
        rom_memory[14470] = 3'b000;
        rom_memory[14471] = 3'b000;
        rom_memory[14472] = 3'b000;
        rom_memory[14473] = 3'b000;
        rom_memory[14474] = 3'b000;
        rom_memory[14475] = 3'b110;
        rom_memory[14476] = 3'b110;
        rom_memory[14477] = 3'b000;
        rom_memory[14478] = 3'b100;
        rom_memory[14479] = 3'b100;
        rom_memory[14480] = 3'b100;
        rom_memory[14481] = 3'b100;
        rom_memory[14482] = 3'b000;
        rom_memory[14483] = 3'b011;
        rom_memory[14484] = 3'b011;
        rom_memory[14485] = 3'b011;
        rom_memory[14486] = 3'b011;
        rom_memory[14487] = 3'b011;
        rom_memory[14488] = 3'b011;
        rom_memory[14489] = 3'b011;
        rom_memory[14490] = 3'b011;
        rom_memory[14491] = 3'b011;
        rom_memory[14492] = 3'b011;
        rom_memory[14493] = 3'b110;
        rom_memory[14494] = 3'b110;
        rom_memory[14495] = 3'b110;
        rom_memory[14496] = 3'b110;
        rom_memory[14497] = 3'b100;
        rom_memory[14498] = 3'b110;
        rom_memory[14499] = 3'b110;
        rom_memory[14500] = 3'b111;
        rom_memory[14501] = 3'b111;
        rom_memory[14502] = 3'b110;
        rom_memory[14503] = 3'b110;
        rom_memory[14504] = 3'b110;
        rom_memory[14505] = 3'b110;
        rom_memory[14506] = 3'b110;
        rom_memory[14507] = 3'b110;
        rom_memory[14508] = 3'b110;
        rom_memory[14509] = 3'b110;
        rom_memory[14510] = 3'b110;
        rom_memory[14511] = 3'b110;
        rom_memory[14512] = 3'b110;
        rom_memory[14513] = 3'b110;
        rom_memory[14514] = 3'b110;
        rom_memory[14515] = 3'b110;
        rom_memory[14516] = 3'b110;
        rom_memory[14517] = 3'b110;
        rom_memory[14518] = 3'b110;
        rom_memory[14519] = 3'b110;
        rom_memory[14520] = 3'b110;
        rom_memory[14521] = 3'b110;
        rom_memory[14522] = 3'b110;
        rom_memory[14523] = 3'b110;
        rom_memory[14524] = 3'b110;
        rom_memory[14525] = 3'b110;
        rom_memory[14526] = 3'b110;
        rom_memory[14527] = 3'b111;
        rom_memory[14528] = 3'b111;
        rom_memory[14529] = 3'b111;
        rom_memory[14530] = 3'b111;
        rom_memory[14531] = 3'b111;
        rom_memory[14532] = 3'b111;
        rom_memory[14533] = 3'b111;
        rom_memory[14534] = 3'b111;
        rom_memory[14535] = 3'b111;
        rom_memory[14536] = 3'b111;
        rom_memory[14537] = 3'b111;
        rom_memory[14538] = 3'b111;
        rom_memory[14539] = 3'b111;
        rom_memory[14540] = 3'b111;
        rom_memory[14541] = 3'b111;
        rom_memory[14542] = 3'b111;
        rom_memory[14543] = 3'b111;
        rom_memory[14544] = 3'b111;
        rom_memory[14545] = 3'b111;
        rom_memory[14546] = 3'b111;
        rom_memory[14547] = 3'b111;
        rom_memory[14548] = 3'b111;
        rom_memory[14549] = 3'b111;
        rom_memory[14550] = 3'b111;
        rom_memory[14551] = 3'b111;
        rom_memory[14552] = 3'b111;
        rom_memory[14553] = 3'b111;
        rom_memory[14554] = 3'b111;
        rom_memory[14555] = 3'b111;
        rom_memory[14556] = 3'b111;
        rom_memory[14557] = 3'b111;
        rom_memory[14558] = 3'b110;
        rom_memory[14559] = 3'b110;
        rom_memory[14560] = 3'b110;
        rom_memory[14561] = 3'b111;
        rom_memory[14562] = 3'b110;
        rom_memory[14563] = 3'b110;
        rom_memory[14564] = 3'b110;
        rom_memory[14565] = 3'b110;
        rom_memory[14566] = 3'b110;
        rom_memory[14567] = 3'b110;
        rom_memory[14568] = 3'b110;
        rom_memory[14569] = 3'b110;
        rom_memory[14570] = 3'b110;
        rom_memory[14571] = 3'b110;
        rom_memory[14572] = 3'b110;
        rom_memory[14573] = 3'b110;
        rom_memory[14574] = 3'b110;
        rom_memory[14575] = 3'b110;
        rom_memory[14576] = 3'b110;
        rom_memory[14577] = 3'b110;
        rom_memory[14578] = 3'b110;
        rom_memory[14579] = 3'b110;
        rom_memory[14580] = 3'b110;
        rom_memory[14581] = 3'b110;
        rom_memory[14582] = 3'b110;
        rom_memory[14583] = 3'b110;
        rom_memory[14584] = 3'b110;
        rom_memory[14585] = 3'b110;
        rom_memory[14586] = 3'b110;
        rom_memory[14587] = 3'b110;
        rom_memory[14588] = 3'b110;
        rom_memory[14589] = 3'b110;
        rom_memory[14590] = 3'b110;
        rom_memory[14591] = 3'b110;
        rom_memory[14592] = 3'b110;
        rom_memory[14593] = 3'b110;
        rom_memory[14594] = 3'b110;
        rom_memory[14595] = 3'b110;
        rom_memory[14596] = 3'b110;
        rom_memory[14597] = 3'b110;
        rom_memory[14598] = 3'b110;
        rom_memory[14599] = 3'b110;
        rom_memory[14600] = 3'b110;
        rom_memory[14601] = 3'b110;
        rom_memory[14602] = 3'b110;
        rom_memory[14603] = 3'b110;
        rom_memory[14604] = 3'b110;
        rom_memory[14605] = 3'b110;
        rom_memory[14606] = 3'b110;
        rom_memory[14607] = 3'b110;
        rom_memory[14608] = 3'b110;
        rom_memory[14609] = 3'b110;
        rom_memory[14610] = 3'b110;
        rom_memory[14611] = 3'b110;
        rom_memory[14612] = 3'b110;
        rom_memory[14613] = 3'b110;
        rom_memory[14614] = 3'b110;
        rom_memory[14615] = 3'b110;
        rom_memory[14616] = 3'b110;
        rom_memory[14617] = 3'b110;
        rom_memory[14618] = 3'b110;
        rom_memory[14619] = 3'b110;
        rom_memory[14620] = 3'b110;
        rom_memory[14621] = 3'b110;
        rom_memory[14622] = 3'b110;
        rom_memory[14623] = 3'b110;
        rom_memory[14624] = 3'b110;
        rom_memory[14625] = 3'b110;
        rom_memory[14626] = 3'b110;
        rom_memory[14627] = 3'b110;
        rom_memory[14628] = 3'b110;
        rom_memory[14629] = 3'b110;
        rom_memory[14630] = 3'b110;
        rom_memory[14631] = 3'b110;
        rom_memory[14632] = 3'b110;
        rom_memory[14633] = 3'b110;
        rom_memory[14634] = 3'b110;
        rom_memory[14635] = 3'b110;
        rom_memory[14636] = 3'b110;
        rom_memory[14637] = 3'b110;
        rom_memory[14638] = 3'b110;
        rom_memory[14639] = 3'b110;
        rom_memory[14640] = 3'b110;
        rom_memory[14641] = 3'b110;
        rom_memory[14642] = 3'b110;
        rom_memory[14643] = 3'b110;
        rom_memory[14644] = 3'b110;
        rom_memory[14645] = 3'b110;
        rom_memory[14646] = 3'b110;
        rom_memory[14647] = 3'b110;
        rom_memory[14648] = 3'b110;
        rom_memory[14649] = 3'b110;
        rom_memory[14650] = 3'b110;
        rom_memory[14651] = 3'b110;
        rom_memory[14652] = 3'b110;
        rom_memory[14653] = 3'b110;
        rom_memory[14654] = 3'b110;
        rom_memory[14655] = 3'b110;
        rom_memory[14656] = 3'b110;
        rom_memory[14657] = 3'b110;
        rom_memory[14658] = 3'b110;
        rom_memory[14659] = 3'b110;
        rom_memory[14660] = 3'b110;
        rom_memory[14661] = 3'b110;
        rom_memory[14662] = 3'b110;
        rom_memory[14663] = 3'b110;
        rom_memory[14664] = 3'b110;
        rom_memory[14665] = 3'b110;
        rom_memory[14666] = 3'b110;
        rom_memory[14667] = 3'b110;
        rom_memory[14668] = 3'b110;
        rom_memory[14669] = 3'b110;
        rom_memory[14670] = 3'b110;
        rom_memory[14671] = 3'b110;
        rom_memory[14672] = 3'b110;
        rom_memory[14673] = 3'b110;
        rom_memory[14674] = 3'b110;
        rom_memory[14675] = 3'b110;
        rom_memory[14676] = 3'b110;
        rom_memory[14677] = 3'b110;
        rom_memory[14678] = 3'b110;
        rom_memory[14679] = 3'b111;
        rom_memory[14680] = 3'b111;
        rom_memory[14681] = 3'b111;
        rom_memory[14682] = 3'b111;
        rom_memory[14683] = 3'b111;
        rom_memory[14684] = 3'b111;
        rom_memory[14685] = 3'b111;
        rom_memory[14686] = 3'b111;
        rom_memory[14687] = 3'b001;
        rom_memory[14688] = 3'b000;
        rom_memory[14689] = 3'b000;
        rom_memory[14690] = 3'b000;
        rom_memory[14691] = 3'b000;
        rom_memory[14692] = 3'b000;
        rom_memory[14693] = 3'b000;
        rom_memory[14694] = 3'b000;
        rom_memory[14695] = 3'b000;
        rom_memory[14696] = 3'b000;
        rom_memory[14697] = 3'b000;
        rom_memory[14698] = 3'b000;
        rom_memory[14699] = 3'b000;
        rom_memory[14700] = 3'b000;
        rom_memory[14701] = 3'b000;
        rom_memory[14702] = 3'b000;
        rom_memory[14703] = 3'b000;
        rom_memory[14704] = 3'b000;
        rom_memory[14705] = 3'b000;
        rom_memory[14706] = 3'b000;
        rom_memory[14707] = 3'b000;
        rom_memory[14708] = 3'b000;
        rom_memory[14709] = 3'b000;
        rom_memory[14710] = 3'b000;
        rom_memory[14711] = 3'b000;
        rom_memory[14712] = 3'b000;
        rom_memory[14713] = 3'b011;
        rom_memory[14714] = 3'b011;
        rom_memory[14715] = 3'b000;
        rom_memory[14716] = 3'b110;
        rom_memory[14717] = 3'b100;
        rom_memory[14718] = 3'b110;
        rom_memory[14719] = 3'b110;
        rom_memory[14720] = 3'b110;
        rom_memory[14721] = 3'b100;
        rom_memory[14722] = 3'b000;
        rom_memory[14723] = 3'b011;
        rom_memory[14724] = 3'b011;
        rom_memory[14725] = 3'b011;
        rom_memory[14726] = 3'b011;
        rom_memory[14727] = 3'b011;
        rom_memory[14728] = 3'b011;
        rom_memory[14729] = 3'b011;
        rom_memory[14730] = 3'b011;
        rom_memory[14731] = 3'b011;
        rom_memory[14732] = 3'b011;
        rom_memory[14733] = 3'b011;
        rom_memory[14734] = 3'b010;
        rom_memory[14735] = 3'b110;
        rom_memory[14736] = 3'b110;
        rom_memory[14737] = 3'b000;
        rom_memory[14738] = 3'b100;
        rom_memory[14739] = 3'b110;
        rom_memory[14740] = 3'b110;
        rom_memory[14741] = 3'b110;
        rom_memory[14742] = 3'b110;
        rom_memory[14743] = 3'b110;
        rom_memory[14744] = 3'b110;
        rom_memory[14745] = 3'b110;
        rom_memory[14746] = 3'b110;
        rom_memory[14747] = 3'b110;
        rom_memory[14748] = 3'b110;
        rom_memory[14749] = 3'b110;
        rom_memory[14750] = 3'b110;
        rom_memory[14751] = 3'b110;
        rom_memory[14752] = 3'b110;
        rom_memory[14753] = 3'b110;
        rom_memory[14754] = 3'b110;
        rom_memory[14755] = 3'b110;
        rom_memory[14756] = 3'b110;
        rom_memory[14757] = 3'b110;
        rom_memory[14758] = 3'b110;
        rom_memory[14759] = 3'b110;
        rom_memory[14760] = 3'b110;
        rom_memory[14761] = 3'b110;
        rom_memory[14762] = 3'b110;
        rom_memory[14763] = 3'b110;
        rom_memory[14764] = 3'b110;
        rom_memory[14765] = 3'b110;
        rom_memory[14766] = 3'b110;
        rom_memory[14767] = 3'b111;
        rom_memory[14768] = 3'b111;
        rom_memory[14769] = 3'b111;
        rom_memory[14770] = 3'b111;
        rom_memory[14771] = 3'b111;
        rom_memory[14772] = 3'b111;
        rom_memory[14773] = 3'b111;
        rom_memory[14774] = 3'b111;
        rom_memory[14775] = 3'b111;
        rom_memory[14776] = 3'b111;
        rom_memory[14777] = 3'b111;
        rom_memory[14778] = 3'b111;
        rom_memory[14779] = 3'b111;
        rom_memory[14780] = 3'b111;
        rom_memory[14781] = 3'b111;
        rom_memory[14782] = 3'b111;
        rom_memory[14783] = 3'b111;
        rom_memory[14784] = 3'b111;
        rom_memory[14785] = 3'b111;
        rom_memory[14786] = 3'b111;
        rom_memory[14787] = 3'b111;
        rom_memory[14788] = 3'b111;
        rom_memory[14789] = 3'b111;
        rom_memory[14790] = 3'b111;
        rom_memory[14791] = 3'b111;
        rom_memory[14792] = 3'b111;
        rom_memory[14793] = 3'b111;
        rom_memory[14794] = 3'b111;
        rom_memory[14795] = 3'b111;
        rom_memory[14796] = 3'b111;
        rom_memory[14797] = 3'b111;
        rom_memory[14798] = 3'b111;
        rom_memory[14799] = 3'b111;
        rom_memory[14800] = 3'b111;
        rom_memory[14801] = 3'b111;
        rom_memory[14802] = 3'b110;
        rom_memory[14803] = 3'b110;
        rom_memory[14804] = 3'b110;
        rom_memory[14805] = 3'b110;
        rom_memory[14806] = 3'b110;
        rom_memory[14807] = 3'b110;
        rom_memory[14808] = 3'b110;
        rom_memory[14809] = 3'b110;
        rom_memory[14810] = 3'b110;
        rom_memory[14811] = 3'b110;
        rom_memory[14812] = 3'b110;
        rom_memory[14813] = 3'b110;
        rom_memory[14814] = 3'b110;
        rom_memory[14815] = 3'b110;
        rom_memory[14816] = 3'b110;
        rom_memory[14817] = 3'b110;
        rom_memory[14818] = 3'b110;
        rom_memory[14819] = 3'b110;
        rom_memory[14820] = 3'b110;
        rom_memory[14821] = 3'b110;
        rom_memory[14822] = 3'b110;
        rom_memory[14823] = 3'b110;
        rom_memory[14824] = 3'b110;
        rom_memory[14825] = 3'b110;
        rom_memory[14826] = 3'b110;
        rom_memory[14827] = 3'b110;
        rom_memory[14828] = 3'b110;
        rom_memory[14829] = 3'b110;
        rom_memory[14830] = 3'b110;
        rom_memory[14831] = 3'b110;
        rom_memory[14832] = 3'b110;
        rom_memory[14833] = 3'b110;
        rom_memory[14834] = 3'b110;
        rom_memory[14835] = 3'b110;
        rom_memory[14836] = 3'b110;
        rom_memory[14837] = 3'b110;
        rom_memory[14838] = 3'b110;
        rom_memory[14839] = 3'b110;
        rom_memory[14840] = 3'b110;
        rom_memory[14841] = 3'b110;
        rom_memory[14842] = 3'b110;
        rom_memory[14843] = 3'b110;
        rom_memory[14844] = 3'b110;
        rom_memory[14845] = 3'b110;
        rom_memory[14846] = 3'b110;
        rom_memory[14847] = 3'b110;
        rom_memory[14848] = 3'b110;
        rom_memory[14849] = 3'b110;
        rom_memory[14850] = 3'b110;
        rom_memory[14851] = 3'b110;
        rom_memory[14852] = 3'b110;
        rom_memory[14853] = 3'b110;
        rom_memory[14854] = 3'b110;
        rom_memory[14855] = 3'b110;
        rom_memory[14856] = 3'b110;
        rom_memory[14857] = 3'b110;
        rom_memory[14858] = 3'b110;
        rom_memory[14859] = 3'b110;
        rom_memory[14860] = 3'b110;
        rom_memory[14861] = 3'b110;
        rom_memory[14862] = 3'b110;
        rom_memory[14863] = 3'b110;
        rom_memory[14864] = 3'b110;
        rom_memory[14865] = 3'b110;
        rom_memory[14866] = 3'b110;
        rom_memory[14867] = 3'b110;
        rom_memory[14868] = 3'b110;
        rom_memory[14869] = 3'b110;
        rom_memory[14870] = 3'b110;
        rom_memory[14871] = 3'b110;
        rom_memory[14872] = 3'b110;
        rom_memory[14873] = 3'b110;
        rom_memory[14874] = 3'b110;
        rom_memory[14875] = 3'b110;
        rom_memory[14876] = 3'b110;
        rom_memory[14877] = 3'b110;
        rom_memory[14878] = 3'b110;
        rom_memory[14879] = 3'b110;
        rom_memory[14880] = 3'b110;
        rom_memory[14881] = 3'b110;
        rom_memory[14882] = 3'b110;
        rom_memory[14883] = 3'b110;
        rom_memory[14884] = 3'b110;
        rom_memory[14885] = 3'b110;
        rom_memory[14886] = 3'b110;
        rom_memory[14887] = 3'b110;
        rom_memory[14888] = 3'b110;
        rom_memory[14889] = 3'b110;
        rom_memory[14890] = 3'b110;
        rom_memory[14891] = 3'b110;
        rom_memory[14892] = 3'b110;
        rom_memory[14893] = 3'b110;
        rom_memory[14894] = 3'b110;
        rom_memory[14895] = 3'b110;
        rom_memory[14896] = 3'b110;
        rom_memory[14897] = 3'b110;
        rom_memory[14898] = 3'b110;
        rom_memory[14899] = 3'b110;
        rom_memory[14900] = 3'b110;
        rom_memory[14901] = 3'b110;
        rom_memory[14902] = 3'b110;
        rom_memory[14903] = 3'b110;
        rom_memory[14904] = 3'b110;
        rom_memory[14905] = 3'b110;
        rom_memory[14906] = 3'b110;
        rom_memory[14907] = 3'b110;
        rom_memory[14908] = 3'b110;
        rom_memory[14909] = 3'b110;
        rom_memory[14910] = 3'b110;
        rom_memory[14911] = 3'b110;
        rom_memory[14912] = 3'b110;
        rom_memory[14913] = 3'b110;
        rom_memory[14914] = 3'b110;
        rom_memory[14915] = 3'b110;
        rom_memory[14916] = 3'b110;
        rom_memory[14917] = 3'b110;
        rom_memory[14918] = 3'b111;
        rom_memory[14919] = 3'b111;
        rom_memory[14920] = 3'b111;
        rom_memory[14921] = 3'b111;
        rom_memory[14922] = 3'b111;
        rom_memory[14923] = 3'b111;
        rom_memory[14924] = 3'b111;
        rom_memory[14925] = 3'b111;
        rom_memory[14926] = 3'b111;
        rom_memory[14927] = 3'b001;
        rom_memory[14928] = 3'b001;
        rom_memory[14929] = 3'b001;
        rom_memory[14930] = 3'b000;
        rom_memory[14931] = 3'b000;
        rom_memory[14932] = 3'b000;
        rom_memory[14933] = 3'b000;
        rom_memory[14934] = 3'b000;
        rom_memory[14935] = 3'b000;
        rom_memory[14936] = 3'b000;
        rom_memory[14937] = 3'b000;
        rom_memory[14938] = 3'b000;
        rom_memory[14939] = 3'b000;
        rom_memory[14940] = 3'b000;
        rom_memory[14941] = 3'b000;
        rom_memory[14942] = 3'b000;
        rom_memory[14943] = 3'b000;
        rom_memory[14944] = 3'b000;
        rom_memory[14945] = 3'b000;
        rom_memory[14946] = 3'b000;
        rom_memory[14947] = 3'b000;
        rom_memory[14948] = 3'b000;
        rom_memory[14949] = 3'b000;
        rom_memory[14950] = 3'b000;
        rom_memory[14951] = 3'b000;
        rom_memory[14952] = 3'b011;
        rom_memory[14953] = 3'b011;
        rom_memory[14954] = 3'b011;
        rom_memory[14955] = 3'b000;
        rom_memory[14956] = 3'b100;
        rom_memory[14957] = 3'b110;
        rom_memory[14958] = 3'b110;
        rom_memory[14959] = 3'b110;
        rom_memory[14960] = 3'b110;
        rom_memory[14961] = 3'b110;
        rom_memory[14962] = 3'b100;
        rom_memory[14963] = 3'b000;
        rom_memory[14964] = 3'b011;
        rom_memory[14965] = 3'b011;
        rom_memory[14966] = 3'b011;
        rom_memory[14967] = 3'b011;
        rom_memory[14968] = 3'b011;
        rom_memory[14969] = 3'b011;
        rom_memory[14970] = 3'b011;
        rom_memory[14971] = 3'b011;
        rom_memory[14972] = 3'b011;
        rom_memory[14973] = 3'b011;
        rom_memory[14974] = 3'b011;
        rom_memory[14975] = 3'b011;
        rom_memory[14976] = 3'b011;
        rom_memory[14977] = 3'b010;
        rom_memory[14978] = 3'b000;
        rom_memory[14979] = 3'b100;
        rom_memory[14980] = 3'b110;
        rom_memory[14981] = 3'b110;
        rom_memory[14982] = 3'b110;
        rom_memory[14983] = 3'b110;
        rom_memory[14984] = 3'b110;
        rom_memory[14985] = 3'b110;
        rom_memory[14986] = 3'b110;
        rom_memory[14987] = 3'b110;
        rom_memory[14988] = 3'b110;
        rom_memory[14989] = 3'b110;
        rom_memory[14990] = 3'b110;
        rom_memory[14991] = 3'b110;
        rom_memory[14992] = 3'b110;
        rom_memory[14993] = 3'b110;
        rom_memory[14994] = 3'b110;
        rom_memory[14995] = 3'b110;
        rom_memory[14996] = 3'b110;
        rom_memory[14997] = 3'b110;
        rom_memory[14998] = 3'b110;
        rom_memory[14999] = 3'b110;
        rom_memory[15000] = 3'b110;
        rom_memory[15001] = 3'b110;
        rom_memory[15002] = 3'b110;
        rom_memory[15003] = 3'b110;
        rom_memory[15004] = 3'b110;
        rom_memory[15005] = 3'b110;
        rom_memory[15006] = 3'b110;
        rom_memory[15007] = 3'b111;
        rom_memory[15008] = 3'b111;
        rom_memory[15009] = 3'b111;
        rom_memory[15010] = 3'b111;
        rom_memory[15011] = 3'b111;
        rom_memory[15012] = 3'b111;
        rom_memory[15013] = 3'b111;
        rom_memory[15014] = 3'b111;
        rom_memory[15015] = 3'b111;
        rom_memory[15016] = 3'b111;
        rom_memory[15017] = 3'b111;
        rom_memory[15018] = 3'b111;
        rom_memory[15019] = 3'b111;
        rom_memory[15020] = 3'b111;
        rom_memory[15021] = 3'b111;
        rom_memory[15022] = 3'b111;
        rom_memory[15023] = 3'b111;
        rom_memory[15024] = 3'b111;
        rom_memory[15025] = 3'b111;
        rom_memory[15026] = 3'b111;
        rom_memory[15027] = 3'b111;
        rom_memory[15028] = 3'b111;
        rom_memory[15029] = 3'b111;
        rom_memory[15030] = 3'b111;
        rom_memory[15031] = 3'b111;
        rom_memory[15032] = 3'b111;
        rom_memory[15033] = 3'b111;
        rom_memory[15034] = 3'b111;
        rom_memory[15035] = 3'b111;
        rom_memory[15036] = 3'b111;
        rom_memory[15037] = 3'b111;
        rom_memory[15038] = 3'b111;
        rom_memory[15039] = 3'b111;
        rom_memory[15040] = 3'b111;
        rom_memory[15041] = 3'b111;
        rom_memory[15042] = 3'b110;
        rom_memory[15043] = 3'b110;
        rom_memory[15044] = 3'b111;
        rom_memory[15045] = 3'b111;
        rom_memory[15046] = 3'b111;
        rom_memory[15047] = 3'b111;
        rom_memory[15048] = 3'b110;
        rom_memory[15049] = 3'b110;
        rom_memory[15050] = 3'b110;
        rom_memory[15051] = 3'b110;
        rom_memory[15052] = 3'b110;
        rom_memory[15053] = 3'b110;
        rom_memory[15054] = 3'b110;
        rom_memory[15055] = 3'b110;
        rom_memory[15056] = 3'b110;
        rom_memory[15057] = 3'b110;
        rom_memory[15058] = 3'b110;
        rom_memory[15059] = 3'b110;
        rom_memory[15060] = 3'b110;
        rom_memory[15061] = 3'b110;
        rom_memory[15062] = 3'b110;
        rom_memory[15063] = 3'b110;
        rom_memory[15064] = 3'b110;
        rom_memory[15065] = 3'b110;
        rom_memory[15066] = 3'b110;
        rom_memory[15067] = 3'b110;
        rom_memory[15068] = 3'b110;
        rom_memory[15069] = 3'b110;
        rom_memory[15070] = 3'b110;
        rom_memory[15071] = 3'b110;
        rom_memory[15072] = 3'b110;
        rom_memory[15073] = 3'b110;
        rom_memory[15074] = 3'b110;
        rom_memory[15075] = 3'b110;
        rom_memory[15076] = 3'b110;
        rom_memory[15077] = 3'b110;
        rom_memory[15078] = 3'b110;
        rom_memory[15079] = 3'b110;
        rom_memory[15080] = 3'b110;
        rom_memory[15081] = 3'b110;
        rom_memory[15082] = 3'b110;
        rom_memory[15083] = 3'b110;
        rom_memory[15084] = 3'b110;
        rom_memory[15085] = 3'b110;
        rom_memory[15086] = 3'b110;
        rom_memory[15087] = 3'b110;
        rom_memory[15088] = 3'b110;
        rom_memory[15089] = 3'b110;
        rom_memory[15090] = 3'b110;
        rom_memory[15091] = 3'b110;
        rom_memory[15092] = 3'b110;
        rom_memory[15093] = 3'b110;
        rom_memory[15094] = 3'b110;
        rom_memory[15095] = 3'b110;
        rom_memory[15096] = 3'b110;
        rom_memory[15097] = 3'b110;
        rom_memory[15098] = 3'b110;
        rom_memory[15099] = 3'b110;
        rom_memory[15100] = 3'b110;
        rom_memory[15101] = 3'b110;
        rom_memory[15102] = 3'b110;
        rom_memory[15103] = 3'b110;
        rom_memory[15104] = 3'b110;
        rom_memory[15105] = 3'b110;
        rom_memory[15106] = 3'b110;
        rom_memory[15107] = 3'b110;
        rom_memory[15108] = 3'b110;
        rom_memory[15109] = 3'b110;
        rom_memory[15110] = 3'b110;
        rom_memory[15111] = 3'b110;
        rom_memory[15112] = 3'b110;
        rom_memory[15113] = 3'b110;
        rom_memory[15114] = 3'b110;
        rom_memory[15115] = 3'b110;
        rom_memory[15116] = 3'b110;
        rom_memory[15117] = 3'b110;
        rom_memory[15118] = 3'b110;
        rom_memory[15119] = 3'b110;
        rom_memory[15120] = 3'b110;
        rom_memory[15121] = 3'b110;
        rom_memory[15122] = 3'b110;
        rom_memory[15123] = 3'b110;
        rom_memory[15124] = 3'b110;
        rom_memory[15125] = 3'b110;
        rom_memory[15126] = 3'b110;
        rom_memory[15127] = 3'b110;
        rom_memory[15128] = 3'b110;
        rom_memory[15129] = 3'b110;
        rom_memory[15130] = 3'b110;
        rom_memory[15131] = 3'b110;
        rom_memory[15132] = 3'b110;
        rom_memory[15133] = 3'b110;
        rom_memory[15134] = 3'b110;
        rom_memory[15135] = 3'b110;
        rom_memory[15136] = 3'b110;
        rom_memory[15137] = 3'b110;
        rom_memory[15138] = 3'b110;
        rom_memory[15139] = 3'b110;
        rom_memory[15140] = 3'b110;
        rom_memory[15141] = 3'b110;
        rom_memory[15142] = 3'b110;
        rom_memory[15143] = 3'b110;
        rom_memory[15144] = 3'b110;
        rom_memory[15145] = 3'b110;
        rom_memory[15146] = 3'b110;
        rom_memory[15147] = 3'b110;
        rom_memory[15148] = 3'b110;
        rom_memory[15149] = 3'b110;
        rom_memory[15150] = 3'b110;
        rom_memory[15151] = 3'b110;
        rom_memory[15152] = 3'b110;
        rom_memory[15153] = 3'b110;
        rom_memory[15154] = 3'b110;
        rom_memory[15155] = 3'b110;
        rom_memory[15156] = 3'b110;
        rom_memory[15157] = 3'b111;
        rom_memory[15158] = 3'b111;
        rom_memory[15159] = 3'b111;
        rom_memory[15160] = 3'b111;
        rom_memory[15161] = 3'b111;
        rom_memory[15162] = 3'b111;
        rom_memory[15163] = 3'b111;
        rom_memory[15164] = 3'b111;
        rom_memory[15165] = 3'b111;
        rom_memory[15166] = 3'b111;
        rom_memory[15167] = 3'b001;
        rom_memory[15168] = 3'b001;
        rom_memory[15169] = 3'b001;
        rom_memory[15170] = 3'b000;
        rom_memory[15171] = 3'b000;
        rom_memory[15172] = 3'b000;
        rom_memory[15173] = 3'b000;
        rom_memory[15174] = 3'b000;
        rom_memory[15175] = 3'b000;
        rom_memory[15176] = 3'b000;
        rom_memory[15177] = 3'b000;
        rom_memory[15178] = 3'b000;
        rom_memory[15179] = 3'b000;
        rom_memory[15180] = 3'b000;
        rom_memory[15181] = 3'b000;
        rom_memory[15182] = 3'b000;
        rom_memory[15183] = 3'b000;
        rom_memory[15184] = 3'b000;
        rom_memory[15185] = 3'b000;
        rom_memory[15186] = 3'b000;
        rom_memory[15187] = 3'b000;
        rom_memory[15188] = 3'b000;
        rom_memory[15189] = 3'b000;
        rom_memory[15190] = 3'b000;
        rom_memory[15191] = 3'b001;
        rom_memory[15192] = 3'b011;
        rom_memory[15193] = 3'b011;
        rom_memory[15194] = 3'b000;
        rom_memory[15195] = 3'b100;
        rom_memory[15196] = 3'b100;
        rom_memory[15197] = 3'b100;
        rom_memory[15198] = 3'b110;
        rom_memory[15199] = 3'b110;
        rom_memory[15200] = 3'b110;
        rom_memory[15201] = 3'b100;
        rom_memory[15202] = 3'b100;
        rom_memory[15203] = 3'b000;
        rom_memory[15204] = 3'b010;
        rom_memory[15205] = 3'b011;
        rom_memory[15206] = 3'b011;
        rom_memory[15207] = 3'b011;
        rom_memory[15208] = 3'b011;
        rom_memory[15209] = 3'b011;
        rom_memory[15210] = 3'b011;
        rom_memory[15211] = 3'b011;
        rom_memory[15212] = 3'b011;
        rom_memory[15213] = 3'b011;
        rom_memory[15214] = 3'b011;
        rom_memory[15215] = 3'b011;
        rom_memory[15216] = 3'b000;
        rom_memory[15217] = 3'b000;
        rom_memory[15218] = 3'b000;
        rom_memory[15219] = 3'b000;
        rom_memory[15220] = 3'b100;
        rom_memory[15221] = 3'b110;
        rom_memory[15222] = 3'b110;
        rom_memory[15223] = 3'b110;
        rom_memory[15224] = 3'b110;
        rom_memory[15225] = 3'b110;
        rom_memory[15226] = 3'b110;
        rom_memory[15227] = 3'b110;
        rom_memory[15228] = 3'b110;
        rom_memory[15229] = 3'b110;
        rom_memory[15230] = 3'b110;
        rom_memory[15231] = 3'b110;
        rom_memory[15232] = 3'b110;
        rom_memory[15233] = 3'b110;
        rom_memory[15234] = 3'b110;
        rom_memory[15235] = 3'b110;
        rom_memory[15236] = 3'b110;
        rom_memory[15237] = 3'b110;
        rom_memory[15238] = 3'b110;
        rom_memory[15239] = 3'b110;
        rom_memory[15240] = 3'b110;
        rom_memory[15241] = 3'b110;
        rom_memory[15242] = 3'b110;
        rom_memory[15243] = 3'b110;
        rom_memory[15244] = 3'b110;
        rom_memory[15245] = 3'b110;
        rom_memory[15246] = 3'b110;
        rom_memory[15247] = 3'b111;
        rom_memory[15248] = 3'b111;
        rom_memory[15249] = 3'b111;
        rom_memory[15250] = 3'b111;
        rom_memory[15251] = 3'b111;
        rom_memory[15252] = 3'b111;
        rom_memory[15253] = 3'b111;
        rom_memory[15254] = 3'b111;
        rom_memory[15255] = 3'b111;
        rom_memory[15256] = 3'b111;
        rom_memory[15257] = 3'b111;
        rom_memory[15258] = 3'b111;
        rom_memory[15259] = 3'b111;
        rom_memory[15260] = 3'b111;
        rom_memory[15261] = 3'b111;
        rom_memory[15262] = 3'b111;
        rom_memory[15263] = 3'b111;
        rom_memory[15264] = 3'b111;
        rom_memory[15265] = 3'b111;
        rom_memory[15266] = 3'b111;
        rom_memory[15267] = 3'b111;
        rom_memory[15268] = 3'b111;
        rom_memory[15269] = 3'b111;
        rom_memory[15270] = 3'b111;
        rom_memory[15271] = 3'b111;
        rom_memory[15272] = 3'b111;
        rom_memory[15273] = 3'b111;
        rom_memory[15274] = 3'b111;
        rom_memory[15275] = 3'b111;
        rom_memory[15276] = 3'b111;
        rom_memory[15277] = 3'b111;
        rom_memory[15278] = 3'b111;
        rom_memory[15279] = 3'b111;
        rom_memory[15280] = 3'b111;
        rom_memory[15281] = 3'b111;
        rom_memory[15282] = 3'b111;
        rom_memory[15283] = 3'b111;
        rom_memory[15284] = 3'b111;
        rom_memory[15285] = 3'b111;
        rom_memory[15286] = 3'b111;
        rom_memory[15287] = 3'b110;
        rom_memory[15288] = 3'b110;
        rom_memory[15289] = 3'b110;
        rom_memory[15290] = 3'b110;
        rom_memory[15291] = 3'b110;
        rom_memory[15292] = 3'b110;
        rom_memory[15293] = 3'b110;
        rom_memory[15294] = 3'b110;
        rom_memory[15295] = 3'b110;
        rom_memory[15296] = 3'b110;
        rom_memory[15297] = 3'b110;
        rom_memory[15298] = 3'b110;
        rom_memory[15299] = 3'b110;
        rom_memory[15300] = 3'b110;
        rom_memory[15301] = 3'b110;
        rom_memory[15302] = 3'b110;
        rom_memory[15303] = 3'b110;
        rom_memory[15304] = 3'b110;
        rom_memory[15305] = 3'b110;
        rom_memory[15306] = 3'b110;
        rom_memory[15307] = 3'b110;
        rom_memory[15308] = 3'b110;
        rom_memory[15309] = 3'b110;
        rom_memory[15310] = 3'b110;
        rom_memory[15311] = 3'b110;
        rom_memory[15312] = 3'b110;
        rom_memory[15313] = 3'b110;
        rom_memory[15314] = 3'b110;
        rom_memory[15315] = 3'b110;
        rom_memory[15316] = 3'b110;
        rom_memory[15317] = 3'b110;
        rom_memory[15318] = 3'b110;
        rom_memory[15319] = 3'b110;
        rom_memory[15320] = 3'b110;
        rom_memory[15321] = 3'b110;
        rom_memory[15322] = 3'b110;
        rom_memory[15323] = 3'b110;
        rom_memory[15324] = 3'b110;
        rom_memory[15325] = 3'b110;
        rom_memory[15326] = 3'b110;
        rom_memory[15327] = 3'b110;
        rom_memory[15328] = 3'b110;
        rom_memory[15329] = 3'b110;
        rom_memory[15330] = 3'b110;
        rom_memory[15331] = 3'b110;
        rom_memory[15332] = 3'b110;
        rom_memory[15333] = 3'b110;
        rom_memory[15334] = 3'b110;
        rom_memory[15335] = 3'b110;
        rom_memory[15336] = 3'b110;
        rom_memory[15337] = 3'b110;
        rom_memory[15338] = 3'b110;
        rom_memory[15339] = 3'b110;
        rom_memory[15340] = 3'b110;
        rom_memory[15341] = 3'b110;
        rom_memory[15342] = 3'b110;
        rom_memory[15343] = 3'b110;
        rom_memory[15344] = 3'b110;
        rom_memory[15345] = 3'b110;
        rom_memory[15346] = 3'b110;
        rom_memory[15347] = 3'b110;
        rom_memory[15348] = 3'b110;
        rom_memory[15349] = 3'b110;
        rom_memory[15350] = 3'b110;
        rom_memory[15351] = 3'b110;
        rom_memory[15352] = 3'b110;
        rom_memory[15353] = 3'b110;
        rom_memory[15354] = 3'b110;
        rom_memory[15355] = 3'b110;
        rom_memory[15356] = 3'b110;
        rom_memory[15357] = 3'b110;
        rom_memory[15358] = 3'b110;
        rom_memory[15359] = 3'b110;
        rom_memory[15360] = 3'b110;
        rom_memory[15361] = 3'b110;
        rom_memory[15362] = 3'b110;
        rom_memory[15363] = 3'b110;
        rom_memory[15364] = 3'b110;
        rom_memory[15365] = 3'b110;
        rom_memory[15366] = 3'b110;
        rom_memory[15367] = 3'b110;
        rom_memory[15368] = 3'b110;
        rom_memory[15369] = 3'b110;
        rom_memory[15370] = 3'b110;
        rom_memory[15371] = 3'b110;
        rom_memory[15372] = 3'b110;
        rom_memory[15373] = 3'b110;
        rom_memory[15374] = 3'b110;
        rom_memory[15375] = 3'b110;
        rom_memory[15376] = 3'b110;
        rom_memory[15377] = 3'b110;
        rom_memory[15378] = 3'b110;
        rom_memory[15379] = 3'b110;
        rom_memory[15380] = 3'b110;
        rom_memory[15381] = 3'b110;
        rom_memory[15382] = 3'b110;
        rom_memory[15383] = 3'b110;
        rom_memory[15384] = 3'b110;
        rom_memory[15385] = 3'b110;
        rom_memory[15386] = 3'b110;
        rom_memory[15387] = 3'b110;
        rom_memory[15388] = 3'b110;
        rom_memory[15389] = 3'b110;
        rom_memory[15390] = 3'b110;
        rom_memory[15391] = 3'b110;
        rom_memory[15392] = 3'b110;
        rom_memory[15393] = 3'b110;
        rom_memory[15394] = 3'b110;
        rom_memory[15395] = 3'b110;
        rom_memory[15396] = 3'b110;
        rom_memory[15397] = 3'b110;
        rom_memory[15398] = 3'b111;
        rom_memory[15399] = 3'b111;
        rom_memory[15400] = 3'b111;
        rom_memory[15401] = 3'b111;
        rom_memory[15402] = 3'b111;
        rom_memory[15403] = 3'b111;
        rom_memory[15404] = 3'b111;
        rom_memory[15405] = 3'b000;
        rom_memory[15406] = 3'b111;
        rom_memory[15407] = 3'b001;
        rom_memory[15408] = 3'b001;
        rom_memory[15409] = 3'b001;
        rom_memory[15410] = 3'b000;
        rom_memory[15411] = 3'b000;
        rom_memory[15412] = 3'b000;
        rom_memory[15413] = 3'b000;
        rom_memory[15414] = 3'b000;
        rom_memory[15415] = 3'b000;
        rom_memory[15416] = 3'b000;
        rom_memory[15417] = 3'b000;
        rom_memory[15418] = 3'b000;
        rom_memory[15419] = 3'b000;
        rom_memory[15420] = 3'b000;
        rom_memory[15421] = 3'b000;
        rom_memory[15422] = 3'b000;
        rom_memory[15423] = 3'b000;
        rom_memory[15424] = 3'b000;
        rom_memory[15425] = 3'b000;
        rom_memory[15426] = 3'b000;
        rom_memory[15427] = 3'b000;
        rom_memory[15428] = 3'b000;
        rom_memory[15429] = 3'b000;
        rom_memory[15430] = 3'b000;
        rom_memory[15431] = 3'b000;
        rom_memory[15432] = 3'b000;
        rom_memory[15433] = 3'b000;
        rom_memory[15434] = 3'b100;
        rom_memory[15435] = 3'b110;
        rom_memory[15436] = 3'b110;
        rom_memory[15437] = 3'b100;
        rom_memory[15438] = 3'b110;
        rom_memory[15439] = 3'b110;
        rom_memory[15440] = 3'b110;
        rom_memory[15441] = 3'b110;
        rom_memory[15442] = 3'b110;
        rom_memory[15443] = 3'b000;
        rom_memory[15444] = 3'b000;
        rom_memory[15445] = 3'b011;
        rom_memory[15446] = 3'b011;
        rom_memory[15447] = 3'b011;
        rom_memory[15448] = 3'b011;
        rom_memory[15449] = 3'b011;
        rom_memory[15450] = 3'b011;
        rom_memory[15451] = 3'b011;
        rom_memory[15452] = 3'b011;
        rom_memory[15453] = 3'b011;
        rom_memory[15454] = 3'b011;
        rom_memory[15455] = 3'b011;
        rom_memory[15456] = 3'b010;
        rom_memory[15457] = 3'b000;
        rom_memory[15458] = 3'b000;
        rom_memory[15459] = 3'b100;
        rom_memory[15460] = 3'b100;
        rom_memory[15461] = 3'b110;
        rom_memory[15462] = 3'b110;
        rom_memory[15463] = 3'b110;
        rom_memory[15464] = 3'b110;
        rom_memory[15465] = 3'b110;
        rom_memory[15466] = 3'b110;
        rom_memory[15467] = 3'b110;
        rom_memory[15468] = 3'b110;
        rom_memory[15469] = 3'b110;
        rom_memory[15470] = 3'b110;
        rom_memory[15471] = 3'b110;
        rom_memory[15472] = 3'b110;
        rom_memory[15473] = 3'b110;
        rom_memory[15474] = 3'b110;
        rom_memory[15475] = 3'b110;
        rom_memory[15476] = 3'b110;
        rom_memory[15477] = 3'b110;
        rom_memory[15478] = 3'b110;
        rom_memory[15479] = 3'b110;
        rom_memory[15480] = 3'b110;
        rom_memory[15481] = 3'b110;
        rom_memory[15482] = 3'b110;
        rom_memory[15483] = 3'b110;
        rom_memory[15484] = 3'b110;
        rom_memory[15485] = 3'b110;
        rom_memory[15486] = 3'b110;
        rom_memory[15487] = 3'b111;
        rom_memory[15488] = 3'b111;
        rom_memory[15489] = 3'b111;
        rom_memory[15490] = 3'b111;
        rom_memory[15491] = 3'b111;
        rom_memory[15492] = 3'b111;
        rom_memory[15493] = 3'b111;
        rom_memory[15494] = 3'b111;
        rom_memory[15495] = 3'b111;
        rom_memory[15496] = 3'b111;
        rom_memory[15497] = 3'b111;
        rom_memory[15498] = 3'b111;
        rom_memory[15499] = 3'b111;
        rom_memory[15500] = 3'b111;
        rom_memory[15501] = 3'b111;
        rom_memory[15502] = 3'b111;
        rom_memory[15503] = 3'b111;
        rom_memory[15504] = 3'b111;
        rom_memory[15505] = 3'b111;
        rom_memory[15506] = 3'b111;
        rom_memory[15507] = 3'b111;
        rom_memory[15508] = 3'b111;
        rom_memory[15509] = 3'b111;
        rom_memory[15510] = 3'b111;
        rom_memory[15511] = 3'b111;
        rom_memory[15512] = 3'b111;
        rom_memory[15513] = 3'b111;
        rom_memory[15514] = 3'b111;
        rom_memory[15515] = 3'b111;
        rom_memory[15516] = 3'b111;
        rom_memory[15517] = 3'b111;
        rom_memory[15518] = 3'b111;
        rom_memory[15519] = 3'b111;
        rom_memory[15520] = 3'b111;
        rom_memory[15521] = 3'b111;
        rom_memory[15522] = 3'b111;
        rom_memory[15523] = 3'b111;
        rom_memory[15524] = 3'b111;
        rom_memory[15525] = 3'b111;
        rom_memory[15526] = 3'b111;
        rom_memory[15527] = 3'b111;
        rom_memory[15528] = 3'b111;
        rom_memory[15529] = 3'b110;
        rom_memory[15530] = 3'b110;
        rom_memory[15531] = 3'b110;
        rom_memory[15532] = 3'b110;
        rom_memory[15533] = 3'b110;
        rom_memory[15534] = 3'b110;
        rom_memory[15535] = 3'b110;
        rom_memory[15536] = 3'b110;
        rom_memory[15537] = 3'b110;
        rom_memory[15538] = 3'b110;
        rom_memory[15539] = 3'b110;
        rom_memory[15540] = 3'b110;
        rom_memory[15541] = 3'b110;
        rom_memory[15542] = 3'b110;
        rom_memory[15543] = 3'b110;
        rom_memory[15544] = 3'b110;
        rom_memory[15545] = 3'b110;
        rom_memory[15546] = 3'b110;
        rom_memory[15547] = 3'b110;
        rom_memory[15548] = 3'b110;
        rom_memory[15549] = 3'b110;
        rom_memory[15550] = 3'b110;
        rom_memory[15551] = 3'b110;
        rom_memory[15552] = 3'b110;
        rom_memory[15553] = 3'b110;
        rom_memory[15554] = 3'b110;
        rom_memory[15555] = 3'b110;
        rom_memory[15556] = 3'b110;
        rom_memory[15557] = 3'b110;
        rom_memory[15558] = 3'b110;
        rom_memory[15559] = 3'b110;
        rom_memory[15560] = 3'b110;
        rom_memory[15561] = 3'b110;
        rom_memory[15562] = 3'b110;
        rom_memory[15563] = 3'b110;
        rom_memory[15564] = 3'b110;
        rom_memory[15565] = 3'b110;
        rom_memory[15566] = 3'b110;
        rom_memory[15567] = 3'b110;
        rom_memory[15568] = 3'b110;
        rom_memory[15569] = 3'b110;
        rom_memory[15570] = 3'b110;
        rom_memory[15571] = 3'b110;
        rom_memory[15572] = 3'b110;
        rom_memory[15573] = 3'b110;
        rom_memory[15574] = 3'b110;
        rom_memory[15575] = 3'b110;
        rom_memory[15576] = 3'b110;
        rom_memory[15577] = 3'b110;
        rom_memory[15578] = 3'b110;
        rom_memory[15579] = 3'b110;
        rom_memory[15580] = 3'b110;
        rom_memory[15581] = 3'b110;
        rom_memory[15582] = 3'b110;
        rom_memory[15583] = 3'b110;
        rom_memory[15584] = 3'b110;
        rom_memory[15585] = 3'b110;
        rom_memory[15586] = 3'b110;
        rom_memory[15587] = 3'b110;
        rom_memory[15588] = 3'b110;
        rom_memory[15589] = 3'b110;
        rom_memory[15590] = 3'b110;
        rom_memory[15591] = 3'b110;
        rom_memory[15592] = 3'b110;
        rom_memory[15593] = 3'b110;
        rom_memory[15594] = 3'b110;
        rom_memory[15595] = 3'b110;
        rom_memory[15596] = 3'b110;
        rom_memory[15597] = 3'b110;
        rom_memory[15598] = 3'b110;
        rom_memory[15599] = 3'b110;
        rom_memory[15600] = 3'b110;
        rom_memory[15601] = 3'b110;
        rom_memory[15602] = 3'b110;
        rom_memory[15603] = 3'b110;
        rom_memory[15604] = 3'b110;
        rom_memory[15605] = 3'b110;
        rom_memory[15606] = 3'b110;
        rom_memory[15607] = 3'b110;
        rom_memory[15608] = 3'b110;
        rom_memory[15609] = 3'b110;
        rom_memory[15610] = 3'b110;
        rom_memory[15611] = 3'b110;
        rom_memory[15612] = 3'b110;
        rom_memory[15613] = 3'b110;
        rom_memory[15614] = 3'b110;
        rom_memory[15615] = 3'b110;
        rom_memory[15616] = 3'b110;
        rom_memory[15617] = 3'b110;
        rom_memory[15618] = 3'b110;
        rom_memory[15619] = 3'b110;
        rom_memory[15620] = 3'b110;
        rom_memory[15621] = 3'b110;
        rom_memory[15622] = 3'b110;
        rom_memory[15623] = 3'b110;
        rom_memory[15624] = 3'b110;
        rom_memory[15625] = 3'b110;
        rom_memory[15626] = 3'b110;
        rom_memory[15627] = 3'b110;
        rom_memory[15628] = 3'b110;
        rom_memory[15629] = 3'b110;
        rom_memory[15630] = 3'b110;
        rom_memory[15631] = 3'b110;
        rom_memory[15632] = 3'b110;
        rom_memory[15633] = 3'b110;
        rom_memory[15634] = 3'b110;
        rom_memory[15635] = 3'b110;
        rom_memory[15636] = 3'b110;
        rom_memory[15637] = 3'b110;
        rom_memory[15638] = 3'b111;
        rom_memory[15639] = 3'b111;
        rom_memory[15640] = 3'b111;
        rom_memory[15641] = 3'b111;
        rom_memory[15642] = 3'b111;
        rom_memory[15643] = 3'b111;
        rom_memory[15644] = 3'b111;
        rom_memory[15645] = 3'b110;
        rom_memory[15646] = 3'b111;
        rom_memory[15647] = 3'b001;
        rom_memory[15648] = 3'b001;
        rom_memory[15649] = 3'b001;
        rom_memory[15650] = 3'b001;
        rom_memory[15651] = 3'b000;
        rom_memory[15652] = 3'b000;
        rom_memory[15653] = 3'b000;
        rom_memory[15654] = 3'b000;
        rom_memory[15655] = 3'b000;
        rom_memory[15656] = 3'b000;
        rom_memory[15657] = 3'b000;
        rom_memory[15658] = 3'b000;
        rom_memory[15659] = 3'b000;
        rom_memory[15660] = 3'b000;
        rom_memory[15661] = 3'b000;
        rom_memory[15662] = 3'b000;
        rom_memory[15663] = 3'b000;
        rom_memory[15664] = 3'b000;
        rom_memory[15665] = 3'b000;
        rom_memory[15666] = 3'b001;
        rom_memory[15667] = 3'b000;
        rom_memory[15668] = 3'b000;
        rom_memory[15669] = 3'b000;
        rom_memory[15670] = 3'b000;
        rom_memory[15671] = 3'b000;
        rom_memory[15672] = 3'b100;
        rom_memory[15673] = 3'b100;
        rom_memory[15674] = 3'b110;
        rom_memory[15675] = 3'b100;
        rom_memory[15676] = 3'b110;
        rom_memory[15677] = 3'b110;
        rom_memory[15678] = 3'b110;
        rom_memory[15679] = 3'b110;
        rom_memory[15680] = 3'b110;
        rom_memory[15681] = 3'b110;
        rom_memory[15682] = 3'b110;
        rom_memory[15683] = 3'b110;
        rom_memory[15684] = 3'b000;
        rom_memory[15685] = 3'b011;
        rom_memory[15686] = 3'b011;
        rom_memory[15687] = 3'b011;
        rom_memory[15688] = 3'b011;
        rom_memory[15689] = 3'b011;
        rom_memory[15690] = 3'b011;
        rom_memory[15691] = 3'b011;
        rom_memory[15692] = 3'b011;
        rom_memory[15693] = 3'b011;
        rom_memory[15694] = 3'b011;
        rom_memory[15695] = 3'b011;
        rom_memory[15696] = 3'b011;
        rom_memory[15697] = 3'b010;
        rom_memory[15698] = 3'b000;
        rom_memory[15699] = 3'b110;
        rom_memory[15700] = 3'b110;
        rom_memory[15701] = 3'b110;
        rom_memory[15702] = 3'b110;
        rom_memory[15703] = 3'b110;
        rom_memory[15704] = 3'b110;
        rom_memory[15705] = 3'b110;
        rom_memory[15706] = 3'b110;
        rom_memory[15707] = 3'b110;
        rom_memory[15708] = 3'b110;
        rom_memory[15709] = 3'b110;
        rom_memory[15710] = 3'b110;
        rom_memory[15711] = 3'b110;
        rom_memory[15712] = 3'b110;
        rom_memory[15713] = 3'b110;
        rom_memory[15714] = 3'b110;
        rom_memory[15715] = 3'b110;
        rom_memory[15716] = 3'b110;
        rom_memory[15717] = 3'b110;
        rom_memory[15718] = 3'b110;
        rom_memory[15719] = 3'b110;
        rom_memory[15720] = 3'b110;
        rom_memory[15721] = 3'b110;
        rom_memory[15722] = 3'b110;
        rom_memory[15723] = 3'b110;
        rom_memory[15724] = 3'b110;
        rom_memory[15725] = 3'b110;
        rom_memory[15726] = 3'b110;
        rom_memory[15727] = 3'b110;
        rom_memory[15728] = 3'b111;
        rom_memory[15729] = 3'b111;
        rom_memory[15730] = 3'b111;
        rom_memory[15731] = 3'b111;
        rom_memory[15732] = 3'b111;
        rom_memory[15733] = 3'b111;
        rom_memory[15734] = 3'b111;
        rom_memory[15735] = 3'b111;
        rom_memory[15736] = 3'b111;
        rom_memory[15737] = 3'b111;
        rom_memory[15738] = 3'b111;
        rom_memory[15739] = 3'b111;
        rom_memory[15740] = 3'b111;
        rom_memory[15741] = 3'b111;
        rom_memory[15742] = 3'b111;
        rom_memory[15743] = 3'b111;
        rom_memory[15744] = 3'b111;
        rom_memory[15745] = 3'b111;
        rom_memory[15746] = 3'b111;
        rom_memory[15747] = 3'b111;
        rom_memory[15748] = 3'b111;
        rom_memory[15749] = 3'b111;
        rom_memory[15750] = 3'b111;
        rom_memory[15751] = 3'b111;
        rom_memory[15752] = 3'b111;
        rom_memory[15753] = 3'b111;
        rom_memory[15754] = 3'b111;
        rom_memory[15755] = 3'b111;
        rom_memory[15756] = 3'b111;
        rom_memory[15757] = 3'b111;
        rom_memory[15758] = 3'b111;
        rom_memory[15759] = 3'b111;
        rom_memory[15760] = 3'b111;
        rom_memory[15761] = 3'b111;
        rom_memory[15762] = 3'b111;
        rom_memory[15763] = 3'b111;
        rom_memory[15764] = 3'b111;
        rom_memory[15765] = 3'b111;
        rom_memory[15766] = 3'b111;
        rom_memory[15767] = 3'b111;
        rom_memory[15768] = 3'b111;
        rom_memory[15769] = 3'b110;
        rom_memory[15770] = 3'b110;
        rom_memory[15771] = 3'b110;
        rom_memory[15772] = 3'b110;
        rom_memory[15773] = 3'b110;
        rom_memory[15774] = 3'b110;
        rom_memory[15775] = 3'b110;
        rom_memory[15776] = 3'b110;
        rom_memory[15777] = 3'b110;
        rom_memory[15778] = 3'b110;
        rom_memory[15779] = 3'b110;
        rom_memory[15780] = 3'b110;
        rom_memory[15781] = 3'b110;
        rom_memory[15782] = 3'b111;
        rom_memory[15783] = 3'b110;
        rom_memory[15784] = 3'b110;
        rom_memory[15785] = 3'b110;
        rom_memory[15786] = 3'b111;
        rom_memory[15787] = 3'b110;
        rom_memory[15788] = 3'b110;
        rom_memory[15789] = 3'b110;
        rom_memory[15790] = 3'b110;
        rom_memory[15791] = 3'b110;
        rom_memory[15792] = 3'b110;
        rom_memory[15793] = 3'b110;
        rom_memory[15794] = 3'b110;
        rom_memory[15795] = 3'b110;
        rom_memory[15796] = 3'b110;
        rom_memory[15797] = 3'b110;
        rom_memory[15798] = 3'b110;
        rom_memory[15799] = 3'b110;
        rom_memory[15800] = 3'b110;
        rom_memory[15801] = 3'b110;
        rom_memory[15802] = 3'b110;
        rom_memory[15803] = 3'b110;
        rom_memory[15804] = 3'b110;
        rom_memory[15805] = 3'b110;
        rom_memory[15806] = 3'b110;
        rom_memory[15807] = 3'b110;
        rom_memory[15808] = 3'b110;
        rom_memory[15809] = 3'b110;
        rom_memory[15810] = 3'b110;
        rom_memory[15811] = 3'b110;
        rom_memory[15812] = 3'b110;
        rom_memory[15813] = 3'b110;
        rom_memory[15814] = 3'b110;
        rom_memory[15815] = 3'b110;
        rom_memory[15816] = 3'b110;
        rom_memory[15817] = 3'b110;
        rom_memory[15818] = 3'b110;
        rom_memory[15819] = 3'b110;
        rom_memory[15820] = 3'b110;
        rom_memory[15821] = 3'b110;
        rom_memory[15822] = 3'b110;
        rom_memory[15823] = 3'b110;
        rom_memory[15824] = 3'b110;
        rom_memory[15825] = 3'b110;
        rom_memory[15826] = 3'b110;
        rom_memory[15827] = 3'b110;
        rom_memory[15828] = 3'b110;
        rom_memory[15829] = 3'b110;
        rom_memory[15830] = 3'b110;
        rom_memory[15831] = 3'b110;
        rom_memory[15832] = 3'b110;
        rom_memory[15833] = 3'b110;
        rom_memory[15834] = 3'b110;
        rom_memory[15835] = 3'b110;
        rom_memory[15836] = 3'b110;
        rom_memory[15837] = 3'b110;
        rom_memory[15838] = 3'b110;
        rom_memory[15839] = 3'b110;
        rom_memory[15840] = 3'b110;
        rom_memory[15841] = 3'b110;
        rom_memory[15842] = 3'b110;
        rom_memory[15843] = 3'b110;
        rom_memory[15844] = 3'b110;
        rom_memory[15845] = 3'b110;
        rom_memory[15846] = 3'b110;
        rom_memory[15847] = 3'b110;
        rom_memory[15848] = 3'b110;
        rom_memory[15849] = 3'b110;
        rom_memory[15850] = 3'b110;
        rom_memory[15851] = 3'b110;
        rom_memory[15852] = 3'b110;
        rom_memory[15853] = 3'b110;
        rom_memory[15854] = 3'b110;
        rom_memory[15855] = 3'b110;
        rom_memory[15856] = 3'b110;
        rom_memory[15857] = 3'b110;
        rom_memory[15858] = 3'b110;
        rom_memory[15859] = 3'b110;
        rom_memory[15860] = 3'b110;
        rom_memory[15861] = 3'b110;
        rom_memory[15862] = 3'b110;
        rom_memory[15863] = 3'b110;
        rom_memory[15864] = 3'b110;
        rom_memory[15865] = 3'b110;
        rom_memory[15866] = 3'b110;
        rom_memory[15867] = 3'b110;
        rom_memory[15868] = 3'b110;
        rom_memory[15869] = 3'b110;
        rom_memory[15870] = 3'b110;
        rom_memory[15871] = 3'b110;
        rom_memory[15872] = 3'b110;
        rom_memory[15873] = 3'b110;
        rom_memory[15874] = 3'b110;
        rom_memory[15875] = 3'b110;
        rom_memory[15876] = 3'b110;
        rom_memory[15877] = 3'b110;
        rom_memory[15878] = 3'b111;
        rom_memory[15879] = 3'b111;
        rom_memory[15880] = 3'b111;
        rom_memory[15881] = 3'b111;
        rom_memory[15882] = 3'b111;
        rom_memory[15883] = 3'b111;
        rom_memory[15884] = 3'b111;
        rom_memory[15885] = 3'b111;
        rom_memory[15886] = 3'b101;
        rom_memory[15887] = 3'b001;
        rom_memory[15888] = 3'b001;
        rom_memory[15889] = 3'b001;
        rom_memory[15890] = 3'b001;
        rom_memory[15891] = 3'b000;
        rom_memory[15892] = 3'b000;
        rom_memory[15893] = 3'b000;
        rom_memory[15894] = 3'b000;
        rom_memory[15895] = 3'b000;
        rom_memory[15896] = 3'b000;
        rom_memory[15897] = 3'b000;
        rom_memory[15898] = 3'b000;
        rom_memory[15899] = 3'b000;
        rom_memory[15900] = 3'b000;
        rom_memory[15901] = 3'b000;
        rom_memory[15902] = 3'b000;
        rom_memory[15903] = 3'b000;
        rom_memory[15904] = 3'b000;
        rom_memory[15905] = 3'b001;
        rom_memory[15906] = 3'b000;
        rom_memory[15907] = 3'b100;
        rom_memory[15908] = 3'b100;
        rom_memory[15909] = 3'b100;
        rom_memory[15910] = 3'b100;
        rom_memory[15911] = 3'b100;
        rom_memory[15912] = 3'b110;
        rom_memory[15913] = 3'b110;
        rom_memory[15914] = 3'b110;
        rom_memory[15915] = 3'b100;
        rom_memory[15916] = 3'b110;
        rom_memory[15917] = 3'b110;
        rom_memory[15918] = 3'b110;
        rom_memory[15919] = 3'b100;
        rom_memory[15920] = 3'b100;
        rom_memory[15921] = 3'b100;
        rom_memory[15922] = 3'b110;
        rom_memory[15923] = 3'b110;
        rom_memory[15924] = 3'b000;
        rom_memory[15925] = 3'b010;
        rom_memory[15926] = 3'b011;
        rom_memory[15927] = 3'b011;
        rom_memory[15928] = 3'b011;
        rom_memory[15929] = 3'b011;
        rom_memory[15930] = 3'b011;
        rom_memory[15931] = 3'b011;
        rom_memory[15932] = 3'b011;
        rom_memory[15933] = 3'b011;
        rom_memory[15934] = 3'b000;
        rom_memory[15935] = 3'b000;
        rom_memory[15936] = 3'b000;
        rom_memory[15937] = 3'b111;
        rom_memory[15938] = 3'b110;
        rom_memory[15939] = 3'b110;
        rom_memory[15940] = 3'b110;
        rom_memory[15941] = 3'b110;
        rom_memory[15942] = 3'b110;
        rom_memory[15943] = 3'b110;
        rom_memory[15944] = 3'b110;
        rom_memory[15945] = 3'b110;
        rom_memory[15946] = 3'b110;
        rom_memory[15947] = 3'b110;
        rom_memory[15948] = 3'b110;
        rom_memory[15949] = 3'b110;
        rom_memory[15950] = 3'b110;
        rom_memory[15951] = 3'b110;
        rom_memory[15952] = 3'b110;
        rom_memory[15953] = 3'b110;
        rom_memory[15954] = 3'b110;
        rom_memory[15955] = 3'b110;
        rom_memory[15956] = 3'b110;
        rom_memory[15957] = 3'b110;
        rom_memory[15958] = 3'b110;
        rom_memory[15959] = 3'b110;
        rom_memory[15960] = 3'b110;
        rom_memory[15961] = 3'b110;
        rom_memory[15962] = 3'b110;
        rom_memory[15963] = 3'b110;
        rom_memory[15964] = 3'b110;
        rom_memory[15965] = 3'b110;
        rom_memory[15966] = 3'b111;
        rom_memory[15967] = 3'b111;
        rom_memory[15968] = 3'b111;
        rom_memory[15969] = 3'b110;
        rom_memory[15970] = 3'b110;
        rom_memory[15971] = 3'b110;
        rom_memory[15972] = 3'b111;
        rom_memory[15973] = 3'b110;
        rom_memory[15974] = 3'b110;
        rom_memory[15975] = 3'b111;
        rom_memory[15976] = 3'b111;
        rom_memory[15977] = 3'b111;
        rom_memory[15978] = 3'b111;
        rom_memory[15979] = 3'b111;
        rom_memory[15980] = 3'b111;
        rom_memory[15981] = 3'b111;
        rom_memory[15982] = 3'b111;
        rom_memory[15983] = 3'b111;
        rom_memory[15984] = 3'b111;
        rom_memory[15985] = 3'b111;
        rom_memory[15986] = 3'b111;
        rom_memory[15987] = 3'b111;
        rom_memory[15988] = 3'b111;
        rom_memory[15989] = 3'b111;
        rom_memory[15990] = 3'b111;
        rom_memory[15991] = 3'b111;
        rom_memory[15992] = 3'b111;
        rom_memory[15993] = 3'b111;
        rom_memory[15994] = 3'b111;
        rom_memory[15995] = 3'b111;
        rom_memory[15996] = 3'b111;
        rom_memory[15997] = 3'b111;
        rom_memory[15998] = 3'b111;
        rom_memory[15999] = 3'b111;
        rom_memory[16000] = 3'b111;
        rom_memory[16001] = 3'b111;
        rom_memory[16002] = 3'b111;
        rom_memory[16003] = 3'b111;
        rom_memory[16004] = 3'b111;
        rom_memory[16005] = 3'b111;
        rom_memory[16006] = 3'b111;
        rom_memory[16007] = 3'b111;
        rom_memory[16008] = 3'b111;
        rom_memory[16009] = 3'b111;
        rom_memory[16010] = 3'b111;
        rom_memory[16011] = 3'b111;
        rom_memory[16012] = 3'b111;
        rom_memory[16013] = 3'b111;
        rom_memory[16014] = 3'b111;
        rom_memory[16015] = 3'b111;
        rom_memory[16016] = 3'b110;
        rom_memory[16017] = 3'b110;
        rom_memory[16018] = 3'b110;
        rom_memory[16019] = 3'b111;
        rom_memory[16020] = 3'b111;
        rom_memory[16021] = 3'b111;
        rom_memory[16022] = 3'b110;
        rom_memory[16023] = 3'b110;
        rom_memory[16024] = 3'b110;
        rom_memory[16025] = 3'b110;
        rom_memory[16026] = 3'b111;
        rom_memory[16027] = 3'b110;
        rom_memory[16028] = 3'b110;
        rom_memory[16029] = 3'b110;
        rom_memory[16030] = 3'b110;
        rom_memory[16031] = 3'b110;
        rom_memory[16032] = 3'b110;
        rom_memory[16033] = 3'b110;
        rom_memory[16034] = 3'b110;
        rom_memory[16035] = 3'b110;
        rom_memory[16036] = 3'b110;
        rom_memory[16037] = 3'b110;
        rom_memory[16038] = 3'b110;
        rom_memory[16039] = 3'b110;
        rom_memory[16040] = 3'b110;
        rom_memory[16041] = 3'b110;
        rom_memory[16042] = 3'b110;
        rom_memory[16043] = 3'b110;
        rom_memory[16044] = 3'b110;
        rom_memory[16045] = 3'b110;
        rom_memory[16046] = 3'b110;
        rom_memory[16047] = 3'b110;
        rom_memory[16048] = 3'b110;
        rom_memory[16049] = 3'b110;
        rom_memory[16050] = 3'b110;
        rom_memory[16051] = 3'b110;
        rom_memory[16052] = 3'b110;
        rom_memory[16053] = 3'b110;
        rom_memory[16054] = 3'b110;
        rom_memory[16055] = 3'b110;
        rom_memory[16056] = 3'b110;
        rom_memory[16057] = 3'b110;
        rom_memory[16058] = 3'b110;
        rom_memory[16059] = 3'b110;
        rom_memory[16060] = 3'b110;
        rom_memory[16061] = 3'b110;
        rom_memory[16062] = 3'b110;
        rom_memory[16063] = 3'b110;
        rom_memory[16064] = 3'b110;
        rom_memory[16065] = 3'b110;
        rom_memory[16066] = 3'b110;
        rom_memory[16067] = 3'b110;
        rom_memory[16068] = 3'b110;
        rom_memory[16069] = 3'b110;
        rom_memory[16070] = 3'b110;
        rom_memory[16071] = 3'b110;
        rom_memory[16072] = 3'b110;
        rom_memory[16073] = 3'b110;
        rom_memory[16074] = 3'b110;
        rom_memory[16075] = 3'b110;
        rom_memory[16076] = 3'b110;
        rom_memory[16077] = 3'b110;
        rom_memory[16078] = 3'b110;
        rom_memory[16079] = 3'b110;
        rom_memory[16080] = 3'b110;
        rom_memory[16081] = 3'b110;
        rom_memory[16082] = 3'b110;
        rom_memory[16083] = 3'b110;
        rom_memory[16084] = 3'b110;
        rom_memory[16085] = 3'b110;
        rom_memory[16086] = 3'b110;
        rom_memory[16087] = 3'b110;
        rom_memory[16088] = 3'b110;
        rom_memory[16089] = 3'b110;
        rom_memory[16090] = 3'b110;
        rom_memory[16091] = 3'b110;
        rom_memory[16092] = 3'b110;
        rom_memory[16093] = 3'b110;
        rom_memory[16094] = 3'b110;
        rom_memory[16095] = 3'b110;
        rom_memory[16096] = 3'b110;
        rom_memory[16097] = 3'b110;
        rom_memory[16098] = 3'b110;
        rom_memory[16099] = 3'b110;
        rom_memory[16100] = 3'b110;
        rom_memory[16101] = 3'b110;
        rom_memory[16102] = 3'b110;
        rom_memory[16103] = 3'b110;
        rom_memory[16104] = 3'b110;
        rom_memory[16105] = 3'b110;
        rom_memory[16106] = 3'b110;
        rom_memory[16107] = 3'b110;
        rom_memory[16108] = 3'b110;
        rom_memory[16109] = 3'b110;
        rom_memory[16110] = 3'b110;
        rom_memory[16111] = 3'b110;
        rom_memory[16112] = 3'b110;
        rom_memory[16113] = 3'b110;
        rom_memory[16114] = 3'b110;
        rom_memory[16115] = 3'b110;
        rom_memory[16116] = 3'b110;
        rom_memory[16117] = 3'b110;
        rom_memory[16118] = 3'b111;
        rom_memory[16119] = 3'b111;
        rom_memory[16120] = 3'b111;
        rom_memory[16121] = 3'b111;
        rom_memory[16122] = 3'b111;
        rom_memory[16123] = 3'b111;
        rom_memory[16124] = 3'b111;
        rom_memory[16125] = 3'b110;
        rom_memory[16126] = 3'b001;
        rom_memory[16127] = 3'b001;
        rom_memory[16128] = 3'b001;
        rom_memory[16129] = 3'b001;
        rom_memory[16130] = 3'b000;
        rom_memory[16131] = 3'b000;
        rom_memory[16132] = 3'b000;
        rom_memory[16133] = 3'b000;
        rom_memory[16134] = 3'b000;
        rom_memory[16135] = 3'b000;
        rom_memory[16136] = 3'b000;
        rom_memory[16137] = 3'b000;
        rom_memory[16138] = 3'b000;
        rom_memory[16139] = 3'b000;
        rom_memory[16140] = 3'b000;
        rom_memory[16141] = 3'b000;
        rom_memory[16142] = 3'b001;
        rom_memory[16143] = 3'b000;
        rom_memory[16144] = 3'b000;
        rom_memory[16145] = 3'b000;
        rom_memory[16146] = 3'b100;
        rom_memory[16147] = 3'b100;
        rom_memory[16148] = 3'b110;
        rom_memory[16149] = 3'b100;
        rom_memory[16150] = 3'b100;
        rom_memory[16151] = 3'b100;
        rom_memory[16152] = 3'b100;
        rom_memory[16153] = 3'b110;
        rom_memory[16154] = 3'b110;
        rom_memory[16155] = 3'b110;
        rom_memory[16156] = 3'b110;
        rom_memory[16157] = 3'b110;
        rom_memory[16158] = 3'b110;
        rom_memory[16159] = 3'b110;
        rom_memory[16160] = 3'b110;
        rom_memory[16161] = 3'b110;
        rom_memory[16162] = 3'b110;
        rom_memory[16163] = 3'b100;
        rom_memory[16164] = 3'b100;
        rom_memory[16165] = 3'b010;
        rom_memory[16166] = 3'b010;
        rom_memory[16167] = 3'b011;
        rom_memory[16168] = 3'b010;
        rom_memory[16169] = 3'b011;
        rom_memory[16170] = 3'b011;
        rom_memory[16171] = 3'b011;
        rom_memory[16172] = 3'b011;
        rom_memory[16173] = 3'b111;
        rom_memory[16174] = 3'b000;
        rom_memory[16175] = 3'b000;
        rom_memory[16176] = 3'b000;
        rom_memory[16177] = 3'b110;
        rom_memory[16178] = 3'b110;
        rom_memory[16179] = 3'b110;
        rom_memory[16180] = 3'b110;
        rom_memory[16181] = 3'b110;
        rom_memory[16182] = 3'b110;
        rom_memory[16183] = 3'b110;
        rom_memory[16184] = 3'b110;
        rom_memory[16185] = 3'b110;
        rom_memory[16186] = 3'b110;
        rom_memory[16187] = 3'b110;
        rom_memory[16188] = 3'b110;
        rom_memory[16189] = 3'b110;
        rom_memory[16190] = 3'b110;
        rom_memory[16191] = 3'b110;
        rom_memory[16192] = 3'b110;
        rom_memory[16193] = 3'b110;
        rom_memory[16194] = 3'b110;
        rom_memory[16195] = 3'b110;
        rom_memory[16196] = 3'b110;
        rom_memory[16197] = 3'b110;
        rom_memory[16198] = 3'b110;
        rom_memory[16199] = 3'b110;
        rom_memory[16200] = 3'b110;
        rom_memory[16201] = 3'b110;
        rom_memory[16202] = 3'b110;
        rom_memory[16203] = 3'b110;
        rom_memory[16204] = 3'b110;
        rom_memory[16205] = 3'b110;
        rom_memory[16206] = 3'b111;
        rom_memory[16207] = 3'b111;
        rom_memory[16208] = 3'b111;
        rom_memory[16209] = 3'b110;
        rom_memory[16210] = 3'b110;
        rom_memory[16211] = 3'b110;
        rom_memory[16212] = 3'b111;
        rom_memory[16213] = 3'b111;
        rom_memory[16214] = 3'b110;
        rom_memory[16215] = 3'b111;
        rom_memory[16216] = 3'b111;
        rom_memory[16217] = 3'b111;
        rom_memory[16218] = 3'b111;
        rom_memory[16219] = 3'b111;
        rom_memory[16220] = 3'b111;
        rom_memory[16221] = 3'b111;
        rom_memory[16222] = 3'b111;
        rom_memory[16223] = 3'b111;
        rom_memory[16224] = 3'b111;
        rom_memory[16225] = 3'b111;
        rom_memory[16226] = 3'b111;
        rom_memory[16227] = 3'b111;
        rom_memory[16228] = 3'b111;
        rom_memory[16229] = 3'b111;
        rom_memory[16230] = 3'b111;
        rom_memory[16231] = 3'b111;
        rom_memory[16232] = 3'b111;
        rom_memory[16233] = 3'b111;
        rom_memory[16234] = 3'b111;
        rom_memory[16235] = 3'b111;
        rom_memory[16236] = 3'b111;
        rom_memory[16237] = 3'b111;
        rom_memory[16238] = 3'b111;
        rom_memory[16239] = 3'b111;
        rom_memory[16240] = 3'b111;
        rom_memory[16241] = 3'b111;
        rom_memory[16242] = 3'b111;
        rom_memory[16243] = 3'b111;
        rom_memory[16244] = 3'b111;
        rom_memory[16245] = 3'b111;
        rom_memory[16246] = 3'b111;
        rom_memory[16247] = 3'b111;
        rom_memory[16248] = 3'b111;
        rom_memory[16249] = 3'b111;
        rom_memory[16250] = 3'b111;
        rom_memory[16251] = 3'b110;
        rom_memory[16252] = 3'b111;
        rom_memory[16253] = 3'b111;
        rom_memory[16254] = 3'b111;
        rom_memory[16255] = 3'b111;
        rom_memory[16256] = 3'b111;
        rom_memory[16257] = 3'b111;
        rom_memory[16258] = 3'b111;
        rom_memory[16259] = 3'b111;
        rom_memory[16260] = 3'b111;
        rom_memory[16261] = 3'b111;
        rom_memory[16262] = 3'b111;
        rom_memory[16263] = 3'b110;
        rom_memory[16264] = 3'b110;
        rom_memory[16265] = 3'b111;
        rom_memory[16266] = 3'b111;
        rom_memory[16267] = 3'b110;
        rom_memory[16268] = 3'b110;
        rom_memory[16269] = 3'b110;
        rom_memory[16270] = 3'b110;
        rom_memory[16271] = 3'b110;
        rom_memory[16272] = 3'b110;
        rom_memory[16273] = 3'b110;
        rom_memory[16274] = 3'b110;
        rom_memory[16275] = 3'b110;
        rom_memory[16276] = 3'b110;
        rom_memory[16277] = 3'b110;
        rom_memory[16278] = 3'b110;
        rom_memory[16279] = 3'b110;
        rom_memory[16280] = 3'b110;
        rom_memory[16281] = 3'b110;
        rom_memory[16282] = 3'b110;
        rom_memory[16283] = 3'b110;
        rom_memory[16284] = 3'b110;
        rom_memory[16285] = 3'b110;
        rom_memory[16286] = 3'b110;
        rom_memory[16287] = 3'b110;
        rom_memory[16288] = 3'b110;
        rom_memory[16289] = 3'b110;
        rom_memory[16290] = 3'b110;
        rom_memory[16291] = 3'b110;
        rom_memory[16292] = 3'b110;
        rom_memory[16293] = 3'b110;
        rom_memory[16294] = 3'b110;
        rom_memory[16295] = 3'b110;
        rom_memory[16296] = 3'b110;
        rom_memory[16297] = 3'b110;
        rom_memory[16298] = 3'b110;
        rom_memory[16299] = 3'b110;
        rom_memory[16300] = 3'b110;
        rom_memory[16301] = 3'b110;
        rom_memory[16302] = 3'b110;
        rom_memory[16303] = 3'b110;
        rom_memory[16304] = 3'b110;
        rom_memory[16305] = 3'b110;
        rom_memory[16306] = 3'b110;
        rom_memory[16307] = 3'b110;
        rom_memory[16308] = 3'b110;
        rom_memory[16309] = 3'b110;
        rom_memory[16310] = 3'b110;
        rom_memory[16311] = 3'b110;
        rom_memory[16312] = 3'b110;
        rom_memory[16313] = 3'b110;
        rom_memory[16314] = 3'b110;
        rom_memory[16315] = 3'b110;
        rom_memory[16316] = 3'b110;
        rom_memory[16317] = 3'b110;
        rom_memory[16318] = 3'b110;
        rom_memory[16319] = 3'b110;
        rom_memory[16320] = 3'b110;
        rom_memory[16321] = 3'b110;
        rom_memory[16322] = 3'b110;
        rom_memory[16323] = 3'b110;
        rom_memory[16324] = 3'b110;
        rom_memory[16325] = 3'b110;
        rom_memory[16326] = 3'b110;
        rom_memory[16327] = 3'b110;
        rom_memory[16328] = 3'b110;
        rom_memory[16329] = 3'b110;
        rom_memory[16330] = 3'b110;
        rom_memory[16331] = 3'b110;
        rom_memory[16332] = 3'b110;
        rom_memory[16333] = 3'b110;
        rom_memory[16334] = 3'b110;
        rom_memory[16335] = 3'b110;
        rom_memory[16336] = 3'b110;
        rom_memory[16337] = 3'b110;
        rom_memory[16338] = 3'b110;
        rom_memory[16339] = 3'b110;
        rom_memory[16340] = 3'b110;
        rom_memory[16341] = 3'b110;
        rom_memory[16342] = 3'b110;
        rom_memory[16343] = 3'b110;
        rom_memory[16344] = 3'b110;
        rom_memory[16345] = 3'b110;
        rom_memory[16346] = 3'b110;
        rom_memory[16347] = 3'b110;
        rom_memory[16348] = 3'b110;
        rom_memory[16349] = 3'b110;
        rom_memory[16350] = 3'b110;
        rom_memory[16351] = 3'b110;
        rom_memory[16352] = 3'b110;
        rom_memory[16353] = 3'b110;
        rom_memory[16354] = 3'b110;
        rom_memory[16355] = 3'b110;
        rom_memory[16356] = 3'b110;
        rom_memory[16357] = 3'b110;
        rom_memory[16358] = 3'b111;
        rom_memory[16359] = 3'b111;
        rom_memory[16360] = 3'b111;
        rom_memory[16361] = 3'b111;
        rom_memory[16362] = 3'b111;
        rom_memory[16363] = 3'b111;
        rom_memory[16364] = 3'b111;
        rom_memory[16365] = 3'b100;
        rom_memory[16366] = 3'b000;
        rom_memory[16367] = 3'b001;
        rom_memory[16368] = 3'b001;
        rom_memory[16369] = 3'b001;
        rom_memory[16370] = 3'b001;
        rom_memory[16371] = 3'b001;
        rom_memory[16372] = 3'b001;
        rom_memory[16373] = 3'b001;
        rom_memory[16374] = 3'b001;
        rom_memory[16375] = 3'b000;
        rom_memory[16376] = 3'b000;
        rom_memory[16377] = 3'b000;
        rom_memory[16378] = 3'b000;
        rom_memory[16379] = 3'b000;
        rom_memory[16380] = 3'b000;
        rom_memory[16381] = 3'b000;
        rom_memory[16382] = 3'b000;
        rom_memory[16383] = 3'b000;
        rom_memory[16384] = 3'b100;
        rom_memory[16385] = 3'b100;
        rom_memory[16386] = 3'b100;
        rom_memory[16387] = 3'b110;
        rom_memory[16388] = 3'b110;
        rom_memory[16389] = 3'b110;
        rom_memory[16390] = 3'b100;
        rom_memory[16391] = 3'b100;
        rom_memory[16392] = 3'b100;
        rom_memory[16393] = 3'b110;
        rom_memory[16394] = 3'b100;
        rom_memory[16395] = 3'b110;
        rom_memory[16396] = 3'b110;
        rom_memory[16397] = 3'b110;
        rom_memory[16398] = 3'b110;
        rom_memory[16399] = 3'b110;
        rom_memory[16400] = 3'b110;
        rom_memory[16401] = 3'b110;
        rom_memory[16402] = 3'b110;
        rom_memory[16403] = 3'b110;
        rom_memory[16404] = 3'b100;
        rom_memory[16405] = 3'b100;
        rom_memory[16406] = 3'b110;
        rom_memory[16407] = 3'b010;
        rom_memory[16408] = 3'b000;
        rom_memory[16409] = 3'b000;
        rom_memory[16410] = 3'b000;
        rom_memory[16411] = 3'b000;
        rom_memory[16412] = 3'b100;
        rom_memory[16413] = 3'b110;
        rom_memory[16414] = 3'b100;
        rom_memory[16415] = 3'b000;
        rom_memory[16416] = 3'b000;
        rom_memory[16417] = 3'b110;
        rom_memory[16418] = 3'b110;
        rom_memory[16419] = 3'b100;
        rom_memory[16420] = 3'b110;
        rom_memory[16421] = 3'b110;
        rom_memory[16422] = 3'b110;
        rom_memory[16423] = 3'b110;
        rom_memory[16424] = 3'b110;
        rom_memory[16425] = 3'b110;
        rom_memory[16426] = 3'b110;
        rom_memory[16427] = 3'b110;
        rom_memory[16428] = 3'b110;
        rom_memory[16429] = 3'b110;
        rom_memory[16430] = 3'b110;
        rom_memory[16431] = 3'b110;
        rom_memory[16432] = 3'b110;
        rom_memory[16433] = 3'b110;
        rom_memory[16434] = 3'b110;
        rom_memory[16435] = 3'b110;
        rom_memory[16436] = 3'b110;
        rom_memory[16437] = 3'b110;
        rom_memory[16438] = 3'b110;
        rom_memory[16439] = 3'b110;
        rom_memory[16440] = 3'b110;
        rom_memory[16441] = 3'b110;
        rom_memory[16442] = 3'b110;
        rom_memory[16443] = 3'b110;
        rom_memory[16444] = 3'b110;
        rom_memory[16445] = 3'b110;
        rom_memory[16446] = 3'b111;
        rom_memory[16447] = 3'b111;
        rom_memory[16448] = 3'b111;
        rom_memory[16449] = 3'b110;
        rom_memory[16450] = 3'b110;
        rom_memory[16451] = 3'b110;
        rom_memory[16452] = 3'b111;
        rom_memory[16453] = 3'b111;
        rom_memory[16454] = 3'b110;
        rom_memory[16455] = 3'b111;
        rom_memory[16456] = 3'b111;
        rom_memory[16457] = 3'b111;
        rom_memory[16458] = 3'b111;
        rom_memory[16459] = 3'b111;
        rom_memory[16460] = 3'b111;
        rom_memory[16461] = 3'b111;
        rom_memory[16462] = 3'b111;
        rom_memory[16463] = 3'b111;
        rom_memory[16464] = 3'b111;
        rom_memory[16465] = 3'b111;
        rom_memory[16466] = 3'b111;
        rom_memory[16467] = 3'b111;
        rom_memory[16468] = 3'b111;
        rom_memory[16469] = 3'b111;
        rom_memory[16470] = 3'b111;
        rom_memory[16471] = 3'b111;
        rom_memory[16472] = 3'b111;
        rom_memory[16473] = 3'b111;
        rom_memory[16474] = 3'b111;
        rom_memory[16475] = 3'b111;
        rom_memory[16476] = 3'b111;
        rom_memory[16477] = 3'b111;
        rom_memory[16478] = 3'b111;
        rom_memory[16479] = 3'b111;
        rom_memory[16480] = 3'b111;
        rom_memory[16481] = 3'b111;
        rom_memory[16482] = 3'b111;
        rom_memory[16483] = 3'b111;
        rom_memory[16484] = 3'b111;
        rom_memory[16485] = 3'b111;
        rom_memory[16486] = 3'b111;
        rom_memory[16487] = 3'b111;
        rom_memory[16488] = 3'b111;
        rom_memory[16489] = 3'b111;
        rom_memory[16490] = 3'b111;
        rom_memory[16491] = 3'b111;
        rom_memory[16492] = 3'b111;
        rom_memory[16493] = 3'b111;
        rom_memory[16494] = 3'b111;
        rom_memory[16495] = 3'b111;
        rom_memory[16496] = 3'b111;
        rom_memory[16497] = 3'b111;
        rom_memory[16498] = 3'b111;
        rom_memory[16499] = 3'b111;
        rom_memory[16500] = 3'b111;
        rom_memory[16501] = 3'b110;
        rom_memory[16502] = 3'b110;
        rom_memory[16503] = 3'b110;
        rom_memory[16504] = 3'b111;
        rom_memory[16505] = 3'b111;
        rom_memory[16506] = 3'b110;
        rom_memory[16507] = 3'b110;
        rom_memory[16508] = 3'b110;
        rom_memory[16509] = 3'b110;
        rom_memory[16510] = 3'b110;
        rom_memory[16511] = 3'b110;
        rom_memory[16512] = 3'b110;
        rom_memory[16513] = 3'b110;
        rom_memory[16514] = 3'b110;
        rom_memory[16515] = 3'b110;
        rom_memory[16516] = 3'b110;
        rom_memory[16517] = 3'b110;
        rom_memory[16518] = 3'b110;
        rom_memory[16519] = 3'b110;
        rom_memory[16520] = 3'b110;
        rom_memory[16521] = 3'b110;
        rom_memory[16522] = 3'b110;
        rom_memory[16523] = 3'b110;
        rom_memory[16524] = 3'b110;
        rom_memory[16525] = 3'b110;
        rom_memory[16526] = 3'b110;
        rom_memory[16527] = 3'b110;
        rom_memory[16528] = 3'b110;
        rom_memory[16529] = 3'b110;
        rom_memory[16530] = 3'b110;
        rom_memory[16531] = 3'b110;
        rom_memory[16532] = 3'b110;
        rom_memory[16533] = 3'b110;
        rom_memory[16534] = 3'b110;
        rom_memory[16535] = 3'b110;
        rom_memory[16536] = 3'b110;
        rom_memory[16537] = 3'b110;
        rom_memory[16538] = 3'b110;
        rom_memory[16539] = 3'b110;
        rom_memory[16540] = 3'b110;
        rom_memory[16541] = 3'b110;
        rom_memory[16542] = 3'b110;
        rom_memory[16543] = 3'b110;
        rom_memory[16544] = 3'b110;
        rom_memory[16545] = 3'b110;
        rom_memory[16546] = 3'b110;
        rom_memory[16547] = 3'b110;
        rom_memory[16548] = 3'b110;
        rom_memory[16549] = 3'b110;
        rom_memory[16550] = 3'b110;
        rom_memory[16551] = 3'b110;
        rom_memory[16552] = 3'b110;
        rom_memory[16553] = 3'b110;
        rom_memory[16554] = 3'b110;
        rom_memory[16555] = 3'b110;
        rom_memory[16556] = 3'b110;
        rom_memory[16557] = 3'b110;
        rom_memory[16558] = 3'b110;
        rom_memory[16559] = 3'b110;
        rom_memory[16560] = 3'b110;
        rom_memory[16561] = 3'b110;
        rom_memory[16562] = 3'b110;
        rom_memory[16563] = 3'b110;
        rom_memory[16564] = 3'b110;
        rom_memory[16565] = 3'b110;
        rom_memory[16566] = 3'b110;
        rom_memory[16567] = 3'b110;
        rom_memory[16568] = 3'b110;
        rom_memory[16569] = 3'b110;
        rom_memory[16570] = 3'b110;
        rom_memory[16571] = 3'b110;
        rom_memory[16572] = 3'b110;
        rom_memory[16573] = 3'b110;
        rom_memory[16574] = 3'b110;
        rom_memory[16575] = 3'b110;
        rom_memory[16576] = 3'b110;
        rom_memory[16577] = 3'b110;
        rom_memory[16578] = 3'b110;
        rom_memory[16579] = 3'b110;
        rom_memory[16580] = 3'b110;
        rom_memory[16581] = 3'b110;
        rom_memory[16582] = 3'b110;
        rom_memory[16583] = 3'b110;
        rom_memory[16584] = 3'b110;
        rom_memory[16585] = 3'b110;
        rom_memory[16586] = 3'b110;
        rom_memory[16587] = 3'b110;
        rom_memory[16588] = 3'b110;
        rom_memory[16589] = 3'b110;
        rom_memory[16590] = 3'b110;
        rom_memory[16591] = 3'b110;
        rom_memory[16592] = 3'b110;
        rom_memory[16593] = 3'b110;
        rom_memory[16594] = 3'b110;
        rom_memory[16595] = 3'b110;
        rom_memory[16596] = 3'b110;
        rom_memory[16597] = 3'b110;
        rom_memory[16598] = 3'b111;
        rom_memory[16599] = 3'b111;
        rom_memory[16600] = 3'b111;
        rom_memory[16601] = 3'b111;
        rom_memory[16602] = 3'b111;
        rom_memory[16603] = 3'b111;
        rom_memory[16604] = 3'b111;
        rom_memory[16605] = 3'b100;
        rom_memory[16606] = 3'b100;
        rom_memory[16607] = 3'b000;
        rom_memory[16608] = 3'b001;
        rom_memory[16609] = 3'b001;
        rom_memory[16610] = 3'b001;
        rom_memory[16611] = 3'b001;
        rom_memory[16612] = 3'b001;
        rom_memory[16613] = 3'b001;
        rom_memory[16614] = 3'b001;
        rom_memory[16615] = 3'b000;
        rom_memory[16616] = 3'b000;
        rom_memory[16617] = 3'b000;
        rom_memory[16618] = 3'b000;
        rom_memory[16619] = 3'b000;
        rom_memory[16620] = 3'b000;
        rom_memory[16621] = 3'b000;
        rom_memory[16622] = 3'b100;
        rom_memory[16623] = 3'b100;
        rom_memory[16624] = 3'b100;
        rom_memory[16625] = 3'b110;
        rom_memory[16626] = 3'b100;
        rom_memory[16627] = 3'b110;
        rom_memory[16628] = 3'b110;
        rom_memory[16629] = 3'b110;
        rom_memory[16630] = 3'b100;
        rom_memory[16631] = 3'b100;
        rom_memory[16632] = 3'b100;
        rom_memory[16633] = 3'b110;
        rom_memory[16634] = 3'b110;
        rom_memory[16635] = 3'b110;
        rom_memory[16636] = 3'b110;
        rom_memory[16637] = 3'b110;
        rom_memory[16638] = 3'b110;
        rom_memory[16639] = 3'b110;
        rom_memory[16640] = 3'b110;
        rom_memory[16641] = 3'b110;
        rom_memory[16642] = 3'b110;
        rom_memory[16643] = 3'b110;
        rom_memory[16644] = 3'b100;
        rom_memory[16645] = 3'b100;
        rom_memory[16646] = 3'b100;
        rom_memory[16647] = 3'b100;
        rom_memory[16648] = 3'b100;
        rom_memory[16649] = 3'b000;
        rom_memory[16650] = 3'b000;
        rom_memory[16651] = 3'b000;
        rom_memory[16652] = 3'b100;
        rom_memory[16653] = 3'b110;
        rom_memory[16654] = 3'b110;
        rom_memory[16655] = 3'b100;
        rom_memory[16656] = 3'b100;
        rom_memory[16657] = 3'b110;
        rom_memory[16658] = 3'b110;
        rom_memory[16659] = 3'b100;
        rom_memory[16660] = 3'b100;
        rom_memory[16661] = 3'b110;
        rom_memory[16662] = 3'b110;
        rom_memory[16663] = 3'b110;
        rom_memory[16664] = 3'b110;
        rom_memory[16665] = 3'b110;
        rom_memory[16666] = 3'b110;
        rom_memory[16667] = 3'b110;
        rom_memory[16668] = 3'b110;
        rom_memory[16669] = 3'b110;
        rom_memory[16670] = 3'b110;
        rom_memory[16671] = 3'b110;
        rom_memory[16672] = 3'b110;
        rom_memory[16673] = 3'b110;
        rom_memory[16674] = 3'b110;
        rom_memory[16675] = 3'b110;
        rom_memory[16676] = 3'b110;
        rom_memory[16677] = 3'b110;
        rom_memory[16678] = 3'b110;
        rom_memory[16679] = 3'b110;
        rom_memory[16680] = 3'b110;
        rom_memory[16681] = 3'b110;
        rom_memory[16682] = 3'b110;
        rom_memory[16683] = 3'b110;
        rom_memory[16684] = 3'b110;
        rom_memory[16685] = 3'b110;
        rom_memory[16686] = 3'b110;
        rom_memory[16687] = 3'b110;
        rom_memory[16688] = 3'b110;
        rom_memory[16689] = 3'b110;
        rom_memory[16690] = 3'b110;
        rom_memory[16691] = 3'b110;
        rom_memory[16692] = 3'b111;
        rom_memory[16693] = 3'b111;
        rom_memory[16694] = 3'b110;
        rom_memory[16695] = 3'b111;
        rom_memory[16696] = 3'b111;
        rom_memory[16697] = 3'b111;
        rom_memory[16698] = 3'b111;
        rom_memory[16699] = 3'b111;
        rom_memory[16700] = 3'b111;
        rom_memory[16701] = 3'b111;
        rom_memory[16702] = 3'b111;
        rom_memory[16703] = 3'b111;
        rom_memory[16704] = 3'b111;
        rom_memory[16705] = 3'b111;
        rom_memory[16706] = 3'b111;
        rom_memory[16707] = 3'b111;
        rom_memory[16708] = 3'b111;
        rom_memory[16709] = 3'b111;
        rom_memory[16710] = 3'b111;
        rom_memory[16711] = 3'b111;
        rom_memory[16712] = 3'b111;
        rom_memory[16713] = 3'b111;
        rom_memory[16714] = 3'b111;
        rom_memory[16715] = 3'b111;
        rom_memory[16716] = 3'b111;
        rom_memory[16717] = 3'b111;
        rom_memory[16718] = 3'b111;
        rom_memory[16719] = 3'b111;
        rom_memory[16720] = 3'b111;
        rom_memory[16721] = 3'b111;
        rom_memory[16722] = 3'b111;
        rom_memory[16723] = 3'b111;
        rom_memory[16724] = 3'b111;
        rom_memory[16725] = 3'b111;
        rom_memory[16726] = 3'b111;
        rom_memory[16727] = 3'b111;
        rom_memory[16728] = 3'b111;
        rom_memory[16729] = 3'b111;
        rom_memory[16730] = 3'b111;
        rom_memory[16731] = 3'b111;
        rom_memory[16732] = 3'b111;
        rom_memory[16733] = 3'b111;
        rom_memory[16734] = 3'b111;
        rom_memory[16735] = 3'b110;
        rom_memory[16736] = 3'b110;
        rom_memory[16737] = 3'b111;
        rom_memory[16738] = 3'b111;
        rom_memory[16739] = 3'b110;
        rom_memory[16740] = 3'b111;
        rom_memory[16741] = 3'b111;
        rom_memory[16742] = 3'b110;
        rom_memory[16743] = 3'b110;
        rom_memory[16744] = 3'b110;
        rom_memory[16745] = 3'b111;
        rom_memory[16746] = 3'b110;
        rom_memory[16747] = 3'b110;
        rom_memory[16748] = 3'b110;
        rom_memory[16749] = 3'b110;
        rom_memory[16750] = 3'b110;
        rom_memory[16751] = 3'b110;
        rom_memory[16752] = 3'b110;
        rom_memory[16753] = 3'b110;
        rom_memory[16754] = 3'b110;
        rom_memory[16755] = 3'b110;
        rom_memory[16756] = 3'b110;
        rom_memory[16757] = 3'b110;
        rom_memory[16758] = 3'b110;
        rom_memory[16759] = 3'b110;
        rom_memory[16760] = 3'b110;
        rom_memory[16761] = 3'b110;
        rom_memory[16762] = 3'b110;
        rom_memory[16763] = 3'b110;
        rom_memory[16764] = 3'b110;
        rom_memory[16765] = 3'b110;
        rom_memory[16766] = 3'b110;
        rom_memory[16767] = 3'b110;
        rom_memory[16768] = 3'b110;
        rom_memory[16769] = 3'b110;
        rom_memory[16770] = 3'b110;
        rom_memory[16771] = 3'b110;
        rom_memory[16772] = 3'b110;
        rom_memory[16773] = 3'b110;
        rom_memory[16774] = 3'b110;
        rom_memory[16775] = 3'b110;
        rom_memory[16776] = 3'b110;
        rom_memory[16777] = 3'b110;
        rom_memory[16778] = 3'b110;
        rom_memory[16779] = 3'b110;
        rom_memory[16780] = 3'b110;
        rom_memory[16781] = 3'b110;
        rom_memory[16782] = 3'b110;
        rom_memory[16783] = 3'b110;
        rom_memory[16784] = 3'b110;
        rom_memory[16785] = 3'b110;
        rom_memory[16786] = 3'b110;
        rom_memory[16787] = 3'b110;
        rom_memory[16788] = 3'b110;
        rom_memory[16789] = 3'b110;
        rom_memory[16790] = 3'b110;
        rom_memory[16791] = 3'b110;
        rom_memory[16792] = 3'b110;
        rom_memory[16793] = 3'b110;
        rom_memory[16794] = 3'b110;
        rom_memory[16795] = 3'b110;
        rom_memory[16796] = 3'b110;
        rom_memory[16797] = 3'b110;
        rom_memory[16798] = 3'b110;
        rom_memory[16799] = 3'b110;
        rom_memory[16800] = 3'b110;
        rom_memory[16801] = 3'b110;
        rom_memory[16802] = 3'b110;
        rom_memory[16803] = 3'b110;
        rom_memory[16804] = 3'b110;
        rom_memory[16805] = 3'b110;
        rom_memory[16806] = 3'b110;
        rom_memory[16807] = 3'b110;
        rom_memory[16808] = 3'b110;
        rom_memory[16809] = 3'b110;
        rom_memory[16810] = 3'b110;
        rom_memory[16811] = 3'b110;
        rom_memory[16812] = 3'b110;
        rom_memory[16813] = 3'b110;
        rom_memory[16814] = 3'b110;
        rom_memory[16815] = 3'b110;
        rom_memory[16816] = 3'b110;
        rom_memory[16817] = 3'b110;
        rom_memory[16818] = 3'b110;
        rom_memory[16819] = 3'b110;
        rom_memory[16820] = 3'b110;
        rom_memory[16821] = 3'b110;
        rom_memory[16822] = 3'b110;
        rom_memory[16823] = 3'b110;
        rom_memory[16824] = 3'b110;
        rom_memory[16825] = 3'b110;
        rom_memory[16826] = 3'b110;
        rom_memory[16827] = 3'b110;
        rom_memory[16828] = 3'b110;
        rom_memory[16829] = 3'b110;
        rom_memory[16830] = 3'b110;
        rom_memory[16831] = 3'b110;
        rom_memory[16832] = 3'b110;
        rom_memory[16833] = 3'b110;
        rom_memory[16834] = 3'b110;
        rom_memory[16835] = 3'b110;
        rom_memory[16836] = 3'b110;
        rom_memory[16837] = 3'b110;
        rom_memory[16838] = 3'b111;
        rom_memory[16839] = 3'b111;
        rom_memory[16840] = 3'b111;
        rom_memory[16841] = 3'b111;
        rom_memory[16842] = 3'b111;
        rom_memory[16843] = 3'b111;
        rom_memory[16844] = 3'b111;
        rom_memory[16845] = 3'b100;
        rom_memory[16846] = 3'b100;
        rom_memory[16847] = 3'b100;
        rom_memory[16848] = 3'b100;
        rom_memory[16849] = 3'b100;
        rom_memory[16850] = 3'b000;
        rom_memory[16851] = 3'b001;
        rom_memory[16852] = 3'b001;
        rom_memory[16853] = 3'b000;
        rom_memory[16854] = 3'b000;
        rom_memory[16855] = 3'b000;
        rom_memory[16856] = 3'b000;
        rom_memory[16857] = 3'b001;
        rom_memory[16858] = 3'b000;
        rom_memory[16859] = 3'b000;
        rom_memory[16860] = 3'b000;
        rom_memory[16861] = 3'b100;
        rom_memory[16862] = 3'b100;
        rom_memory[16863] = 3'b100;
        rom_memory[16864] = 3'b100;
        rom_memory[16865] = 3'b110;
        rom_memory[16866] = 3'b100;
        rom_memory[16867] = 3'b100;
        rom_memory[16868] = 3'b110;
        rom_memory[16869] = 3'b110;
        rom_memory[16870] = 3'b100;
        rom_memory[16871] = 3'b100;
        rom_memory[16872] = 3'b100;
        rom_memory[16873] = 3'b100;
        rom_memory[16874] = 3'b110;
        rom_memory[16875] = 3'b110;
        rom_memory[16876] = 3'b110;
        rom_memory[16877] = 3'b110;
        rom_memory[16878] = 3'b110;
        rom_memory[16879] = 3'b110;
        rom_memory[16880] = 3'b110;
        rom_memory[16881] = 3'b110;
        rom_memory[16882] = 3'b110;
        rom_memory[16883] = 3'b110;
        rom_memory[16884] = 3'b110;
        rom_memory[16885] = 3'b100;
        rom_memory[16886] = 3'b000;
        rom_memory[16887] = 3'b100;
        rom_memory[16888] = 3'b100;
        rom_memory[16889] = 3'b100;
        rom_memory[16890] = 3'b100;
        rom_memory[16891] = 3'b000;
        rom_memory[16892] = 3'b000;
        rom_memory[16893] = 3'b110;
        rom_memory[16894] = 3'b110;
        rom_memory[16895] = 3'b110;
        rom_memory[16896] = 3'b110;
        rom_memory[16897] = 3'b110;
        rom_memory[16898] = 3'b110;
        rom_memory[16899] = 3'b110;
        rom_memory[16900] = 3'b110;
        rom_memory[16901] = 3'b110;
        rom_memory[16902] = 3'b110;
        rom_memory[16903] = 3'b110;
        rom_memory[16904] = 3'b110;
        rom_memory[16905] = 3'b110;
        rom_memory[16906] = 3'b110;
        rom_memory[16907] = 3'b110;
        rom_memory[16908] = 3'b110;
        rom_memory[16909] = 3'b110;
        rom_memory[16910] = 3'b110;
        rom_memory[16911] = 3'b110;
        rom_memory[16912] = 3'b110;
        rom_memory[16913] = 3'b110;
        rom_memory[16914] = 3'b110;
        rom_memory[16915] = 3'b110;
        rom_memory[16916] = 3'b110;
        rom_memory[16917] = 3'b110;
        rom_memory[16918] = 3'b110;
        rom_memory[16919] = 3'b110;
        rom_memory[16920] = 3'b110;
        rom_memory[16921] = 3'b110;
        rom_memory[16922] = 3'b110;
        rom_memory[16923] = 3'b110;
        rom_memory[16924] = 3'b110;
        rom_memory[16925] = 3'b110;
        rom_memory[16926] = 3'b110;
        rom_memory[16927] = 3'b110;
        rom_memory[16928] = 3'b110;
        rom_memory[16929] = 3'b111;
        rom_memory[16930] = 3'b110;
        rom_memory[16931] = 3'b110;
        rom_memory[16932] = 3'b111;
        rom_memory[16933] = 3'b110;
        rom_memory[16934] = 3'b111;
        rom_memory[16935] = 3'b111;
        rom_memory[16936] = 3'b111;
        rom_memory[16937] = 3'b111;
        rom_memory[16938] = 3'b111;
        rom_memory[16939] = 3'b111;
        rom_memory[16940] = 3'b111;
        rom_memory[16941] = 3'b111;
        rom_memory[16942] = 3'b111;
        rom_memory[16943] = 3'b111;
        rom_memory[16944] = 3'b111;
        rom_memory[16945] = 3'b111;
        rom_memory[16946] = 3'b111;
        rom_memory[16947] = 3'b111;
        rom_memory[16948] = 3'b111;
        rom_memory[16949] = 3'b111;
        rom_memory[16950] = 3'b111;
        rom_memory[16951] = 3'b111;
        rom_memory[16952] = 3'b111;
        rom_memory[16953] = 3'b111;
        rom_memory[16954] = 3'b111;
        rom_memory[16955] = 3'b111;
        rom_memory[16956] = 3'b111;
        rom_memory[16957] = 3'b111;
        rom_memory[16958] = 3'b111;
        rom_memory[16959] = 3'b111;
        rom_memory[16960] = 3'b111;
        rom_memory[16961] = 3'b111;
        rom_memory[16962] = 3'b111;
        rom_memory[16963] = 3'b111;
        rom_memory[16964] = 3'b111;
        rom_memory[16965] = 3'b111;
        rom_memory[16966] = 3'b111;
        rom_memory[16967] = 3'b111;
        rom_memory[16968] = 3'b111;
        rom_memory[16969] = 3'b111;
        rom_memory[16970] = 3'b111;
        rom_memory[16971] = 3'b111;
        rom_memory[16972] = 3'b111;
        rom_memory[16973] = 3'b111;
        rom_memory[16974] = 3'b111;
        rom_memory[16975] = 3'b111;
        rom_memory[16976] = 3'b111;
        rom_memory[16977] = 3'b110;
        rom_memory[16978] = 3'b111;
        rom_memory[16979] = 3'b111;
        rom_memory[16980] = 3'b111;
        rom_memory[16981] = 3'b111;
        rom_memory[16982] = 3'b110;
        rom_memory[16983] = 3'b110;
        rom_memory[16984] = 3'b110;
        rom_memory[16985] = 3'b111;
        rom_memory[16986] = 3'b110;
        rom_memory[16987] = 3'b110;
        rom_memory[16988] = 3'b110;
        rom_memory[16989] = 3'b111;
        rom_memory[16990] = 3'b110;
        rom_memory[16991] = 3'b110;
        rom_memory[16992] = 3'b110;
        rom_memory[16993] = 3'b110;
        rom_memory[16994] = 3'b110;
        rom_memory[16995] = 3'b110;
        rom_memory[16996] = 3'b110;
        rom_memory[16997] = 3'b110;
        rom_memory[16998] = 3'b110;
        rom_memory[16999] = 3'b110;
        rom_memory[17000] = 3'b110;
        rom_memory[17001] = 3'b110;
        rom_memory[17002] = 3'b110;
        rom_memory[17003] = 3'b110;
        rom_memory[17004] = 3'b110;
        rom_memory[17005] = 3'b110;
        rom_memory[17006] = 3'b110;
        rom_memory[17007] = 3'b110;
        rom_memory[17008] = 3'b110;
        rom_memory[17009] = 3'b110;
        rom_memory[17010] = 3'b110;
        rom_memory[17011] = 3'b110;
        rom_memory[17012] = 3'b110;
        rom_memory[17013] = 3'b110;
        rom_memory[17014] = 3'b110;
        rom_memory[17015] = 3'b110;
        rom_memory[17016] = 3'b110;
        rom_memory[17017] = 3'b110;
        rom_memory[17018] = 3'b110;
        rom_memory[17019] = 3'b110;
        rom_memory[17020] = 3'b110;
        rom_memory[17021] = 3'b110;
        rom_memory[17022] = 3'b110;
        rom_memory[17023] = 3'b110;
        rom_memory[17024] = 3'b110;
        rom_memory[17025] = 3'b110;
        rom_memory[17026] = 3'b110;
        rom_memory[17027] = 3'b110;
        rom_memory[17028] = 3'b110;
        rom_memory[17029] = 3'b110;
        rom_memory[17030] = 3'b110;
        rom_memory[17031] = 3'b110;
        rom_memory[17032] = 3'b110;
        rom_memory[17033] = 3'b110;
        rom_memory[17034] = 3'b110;
        rom_memory[17035] = 3'b110;
        rom_memory[17036] = 3'b110;
        rom_memory[17037] = 3'b110;
        rom_memory[17038] = 3'b110;
        rom_memory[17039] = 3'b110;
        rom_memory[17040] = 3'b110;
        rom_memory[17041] = 3'b110;
        rom_memory[17042] = 3'b110;
        rom_memory[17043] = 3'b110;
        rom_memory[17044] = 3'b110;
        rom_memory[17045] = 3'b110;
        rom_memory[17046] = 3'b110;
        rom_memory[17047] = 3'b110;
        rom_memory[17048] = 3'b110;
        rom_memory[17049] = 3'b110;
        rom_memory[17050] = 3'b110;
        rom_memory[17051] = 3'b110;
        rom_memory[17052] = 3'b110;
        rom_memory[17053] = 3'b110;
        rom_memory[17054] = 3'b110;
        rom_memory[17055] = 3'b110;
        rom_memory[17056] = 3'b110;
        rom_memory[17057] = 3'b110;
        rom_memory[17058] = 3'b110;
        rom_memory[17059] = 3'b110;
        rom_memory[17060] = 3'b110;
        rom_memory[17061] = 3'b110;
        rom_memory[17062] = 3'b110;
        rom_memory[17063] = 3'b110;
        rom_memory[17064] = 3'b110;
        rom_memory[17065] = 3'b110;
        rom_memory[17066] = 3'b110;
        rom_memory[17067] = 3'b110;
        rom_memory[17068] = 3'b110;
        rom_memory[17069] = 3'b110;
        rom_memory[17070] = 3'b110;
        rom_memory[17071] = 3'b110;
        rom_memory[17072] = 3'b110;
        rom_memory[17073] = 3'b110;
        rom_memory[17074] = 3'b110;
        rom_memory[17075] = 3'b110;
        rom_memory[17076] = 3'b111;
        rom_memory[17077] = 3'b111;
        rom_memory[17078] = 3'b111;
        rom_memory[17079] = 3'b111;
        rom_memory[17080] = 3'b111;
        rom_memory[17081] = 3'b111;
        rom_memory[17082] = 3'b111;
        rom_memory[17083] = 3'b111;
        rom_memory[17084] = 3'b111;
        rom_memory[17085] = 3'b110;
        rom_memory[17086] = 3'b100;
        rom_memory[17087] = 3'b100;
        rom_memory[17088] = 3'b100;
        rom_memory[17089] = 3'b100;
        rom_memory[17090] = 3'b100;
        rom_memory[17091] = 3'b000;
        rom_memory[17092] = 3'b000;
        rom_memory[17093] = 3'b000;
        rom_memory[17094] = 3'b000;
        rom_memory[17095] = 3'b000;
        rom_memory[17096] = 3'b000;
        rom_memory[17097] = 3'b000;
        rom_memory[17098] = 3'b000;
        rom_memory[17099] = 3'b000;
        rom_memory[17100] = 3'b100;
        rom_memory[17101] = 3'b100;
        rom_memory[17102] = 3'b100;
        rom_memory[17103] = 3'b100;
        rom_memory[17104] = 3'b100;
        rom_memory[17105] = 3'b100;
        rom_memory[17106] = 3'b110;
        rom_memory[17107] = 3'b100;
        rom_memory[17108] = 3'b110;
        rom_memory[17109] = 3'b110;
        rom_memory[17110] = 3'b100;
        rom_memory[17111] = 3'b100;
        rom_memory[17112] = 3'b110;
        rom_memory[17113] = 3'b100;
        rom_memory[17114] = 3'b110;
        rom_memory[17115] = 3'b110;
        rom_memory[17116] = 3'b110;
        rom_memory[17117] = 3'b110;
        rom_memory[17118] = 3'b110;
        rom_memory[17119] = 3'b110;
        rom_memory[17120] = 3'b110;
        rom_memory[17121] = 3'b110;
        rom_memory[17122] = 3'b110;
        rom_memory[17123] = 3'b110;
        rom_memory[17124] = 3'b110;
        rom_memory[17125] = 3'b110;
        rom_memory[17126] = 3'b110;
        rom_memory[17127] = 3'b100;
        rom_memory[17128] = 3'b100;
        rom_memory[17129] = 3'b100;
        rom_memory[17130] = 3'b100;
        rom_memory[17131] = 3'b000;
        rom_memory[17132] = 3'b000;
        rom_memory[17133] = 3'b100;
        rom_memory[17134] = 3'b100;
        rom_memory[17135] = 3'b110;
        rom_memory[17136] = 3'b110;
        rom_memory[17137] = 3'b110;
        rom_memory[17138] = 3'b110;
        rom_memory[17139] = 3'b110;
        rom_memory[17140] = 3'b110;
        rom_memory[17141] = 3'b111;
        rom_memory[17142] = 3'b110;
        rom_memory[17143] = 3'b100;
        rom_memory[17144] = 3'b110;
        rom_memory[17145] = 3'b110;
        rom_memory[17146] = 3'b110;
        rom_memory[17147] = 3'b110;
        rom_memory[17148] = 3'b110;
        rom_memory[17149] = 3'b111;
        rom_memory[17150] = 3'b111;
        rom_memory[17151] = 3'b111;
        rom_memory[17152] = 3'b110;
        rom_memory[17153] = 3'b110;
        rom_memory[17154] = 3'b110;
        rom_memory[17155] = 3'b110;
        rom_memory[17156] = 3'b110;
        rom_memory[17157] = 3'b110;
        rom_memory[17158] = 3'b110;
        rom_memory[17159] = 3'b110;
        rom_memory[17160] = 3'b110;
        rom_memory[17161] = 3'b110;
        rom_memory[17162] = 3'b110;
        rom_memory[17163] = 3'b110;
        rom_memory[17164] = 3'b110;
        rom_memory[17165] = 3'b110;
        rom_memory[17166] = 3'b111;
        rom_memory[17167] = 3'b111;
        rom_memory[17168] = 3'b111;
        rom_memory[17169] = 3'b110;
        rom_memory[17170] = 3'b111;
        rom_memory[17171] = 3'b111;
        rom_memory[17172] = 3'b111;
        rom_memory[17173] = 3'b110;
        rom_memory[17174] = 3'b110;
        rom_memory[17175] = 3'b111;
        rom_memory[17176] = 3'b111;
        rom_memory[17177] = 3'b111;
        rom_memory[17178] = 3'b111;
        rom_memory[17179] = 3'b111;
        rom_memory[17180] = 3'b111;
        rom_memory[17181] = 3'b111;
        rom_memory[17182] = 3'b111;
        rom_memory[17183] = 3'b111;
        rom_memory[17184] = 3'b111;
        rom_memory[17185] = 3'b111;
        rom_memory[17186] = 3'b111;
        rom_memory[17187] = 3'b111;
        rom_memory[17188] = 3'b111;
        rom_memory[17189] = 3'b111;
        rom_memory[17190] = 3'b111;
        rom_memory[17191] = 3'b111;
        rom_memory[17192] = 3'b111;
        rom_memory[17193] = 3'b111;
        rom_memory[17194] = 3'b111;
        rom_memory[17195] = 3'b111;
        rom_memory[17196] = 3'b111;
        rom_memory[17197] = 3'b111;
        rom_memory[17198] = 3'b111;
        rom_memory[17199] = 3'b111;
        rom_memory[17200] = 3'b111;
        rom_memory[17201] = 3'b111;
        rom_memory[17202] = 3'b111;
        rom_memory[17203] = 3'b111;
        rom_memory[17204] = 3'b111;
        rom_memory[17205] = 3'b111;
        rom_memory[17206] = 3'b111;
        rom_memory[17207] = 3'b111;
        rom_memory[17208] = 3'b111;
        rom_memory[17209] = 3'b111;
        rom_memory[17210] = 3'b111;
        rom_memory[17211] = 3'b111;
        rom_memory[17212] = 3'b111;
        rom_memory[17213] = 3'b111;
        rom_memory[17214] = 3'b111;
        rom_memory[17215] = 3'b111;
        rom_memory[17216] = 3'b111;
        rom_memory[17217] = 3'b111;
        rom_memory[17218] = 3'b111;
        rom_memory[17219] = 3'b111;
        rom_memory[17220] = 3'b111;
        rom_memory[17221] = 3'b111;
        rom_memory[17222] = 3'b111;
        rom_memory[17223] = 3'b110;
        rom_memory[17224] = 3'b110;
        rom_memory[17225] = 3'b111;
        rom_memory[17226] = 3'b110;
        rom_memory[17227] = 3'b110;
        rom_memory[17228] = 3'b111;
        rom_memory[17229] = 3'b111;
        rom_memory[17230] = 3'b110;
        rom_memory[17231] = 3'b110;
        rom_memory[17232] = 3'b110;
        rom_memory[17233] = 3'b110;
        rom_memory[17234] = 3'b110;
        rom_memory[17235] = 3'b110;
        rom_memory[17236] = 3'b110;
        rom_memory[17237] = 3'b110;
        rom_memory[17238] = 3'b110;
        rom_memory[17239] = 3'b110;
        rom_memory[17240] = 3'b110;
        rom_memory[17241] = 3'b110;
        rom_memory[17242] = 3'b110;
        rom_memory[17243] = 3'b110;
        rom_memory[17244] = 3'b110;
        rom_memory[17245] = 3'b110;
        rom_memory[17246] = 3'b110;
        rom_memory[17247] = 3'b110;
        rom_memory[17248] = 3'b110;
        rom_memory[17249] = 3'b110;
        rom_memory[17250] = 3'b110;
        rom_memory[17251] = 3'b110;
        rom_memory[17252] = 3'b110;
        rom_memory[17253] = 3'b110;
        rom_memory[17254] = 3'b110;
        rom_memory[17255] = 3'b110;
        rom_memory[17256] = 3'b110;
        rom_memory[17257] = 3'b110;
        rom_memory[17258] = 3'b110;
        rom_memory[17259] = 3'b110;
        rom_memory[17260] = 3'b110;
        rom_memory[17261] = 3'b110;
        rom_memory[17262] = 3'b110;
        rom_memory[17263] = 3'b110;
        rom_memory[17264] = 3'b110;
        rom_memory[17265] = 3'b110;
        rom_memory[17266] = 3'b110;
        rom_memory[17267] = 3'b110;
        rom_memory[17268] = 3'b110;
        rom_memory[17269] = 3'b110;
        rom_memory[17270] = 3'b110;
        rom_memory[17271] = 3'b110;
        rom_memory[17272] = 3'b110;
        rom_memory[17273] = 3'b110;
        rom_memory[17274] = 3'b110;
        rom_memory[17275] = 3'b110;
        rom_memory[17276] = 3'b110;
        rom_memory[17277] = 3'b110;
        rom_memory[17278] = 3'b110;
        rom_memory[17279] = 3'b110;
        rom_memory[17280] = 3'b110;
        rom_memory[17281] = 3'b110;
        rom_memory[17282] = 3'b110;
        rom_memory[17283] = 3'b110;
        rom_memory[17284] = 3'b110;
        rom_memory[17285] = 3'b110;
        rom_memory[17286] = 3'b110;
        rom_memory[17287] = 3'b110;
        rom_memory[17288] = 3'b110;
        rom_memory[17289] = 3'b110;
        rom_memory[17290] = 3'b110;
        rom_memory[17291] = 3'b110;
        rom_memory[17292] = 3'b110;
        rom_memory[17293] = 3'b110;
        rom_memory[17294] = 3'b110;
        rom_memory[17295] = 3'b110;
        rom_memory[17296] = 3'b110;
        rom_memory[17297] = 3'b110;
        rom_memory[17298] = 3'b110;
        rom_memory[17299] = 3'b110;
        rom_memory[17300] = 3'b110;
        rom_memory[17301] = 3'b110;
        rom_memory[17302] = 3'b110;
        rom_memory[17303] = 3'b110;
        rom_memory[17304] = 3'b110;
        rom_memory[17305] = 3'b110;
        rom_memory[17306] = 3'b110;
        rom_memory[17307] = 3'b110;
        rom_memory[17308] = 3'b110;
        rom_memory[17309] = 3'b110;
        rom_memory[17310] = 3'b110;
        rom_memory[17311] = 3'b110;
        rom_memory[17312] = 3'b110;
        rom_memory[17313] = 3'b110;
        rom_memory[17314] = 3'b110;
        rom_memory[17315] = 3'b110;
        rom_memory[17316] = 3'b111;
        rom_memory[17317] = 3'b111;
        rom_memory[17318] = 3'b111;
        rom_memory[17319] = 3'b111;
        rom_memory[17320] = 3'b111;
        rom_memory[17321] = 3'b111;
        rom_memory[17322] = 3'b111;
        rom_memory[17323] = 3'b111;
        rom_memory[17324] = 3'b111;
        rom_memory[17325] = 3'b110;
        rom_memory[17326] = 3'b100;
        rom_memory[17327] = 3'b100;
        rom_memory[17328] = 3'b100;
        rom_memory[17329] = 3'b100;
        rom_memory[17330] = 3'b100;
        rom_memory[17331] = 3'b100;
        rom_memory[17332] = 3'b100;
        rom_memory[17333] = 3'b100;
        rom_memory[17334] = 3'b100;
        rom_memory[17335] = 3'b100;
        rom_memory[17336] = 3'b000;
        rom_memory[17337] = 3'b000;
        rom_memory[17338] = 3'b000;
        rom_memory[17339] = 3'b100;
        rom_memory[17340] = 3'b100;
        rom_memory[17341] = 3'b100;
        rom_memory[17342] = 3'b100;
        rom_memory[17343] = 3'b100;
        rom_memory[17344] = 3'b110;
        rom_memory[17345] = 3'b110;
        rom_memory[17346] = 3'b110;
        rom_memory[17347] = 3'b110;
        rom_memory[17348] = 3'b100;
        rom_memory[17349] = 3'b110;
        rom_memory[17350] = 3'b100;
        rom_memory[17351] = 3'b100;
        rom_memory[17352] = 3'b110;
        rom_memory[17353] = 3'b110;
        rom_memory[17354] = 3'b110;
        rom_memory[17355] = 3'b110;
        rom_memory[17356] = 3'b110;
        rom_memory[17357] = 3'b110;
        rom_memory[17358] = 3'b110;
        rom_memory[17359] = 3'b110;
        rom_memory[17360] = 3'b110;
        rom_memory[17361] = 3'b110;
        rom_memory[17362] = 3'b110;
        rom_memory[17363] = 3'b110;
        rom_memory[17364] = 3'b110;
        rom_memory[17365] = 3'b110;
        rom_memory[17366] = 3'b110;
        rom_memory[17367] = 3'b110;
        rom_memory[17368] = 3'b110;
        rom_memory[17369] = 3'b100;
        rom_memory[17370] = 3'b000;
        rom_memory[17371] = 3'b000;
        rom_memory[17372] = 3'b000;
        rom_memory[17373] = 3'b000;
        rom_memory[17374] = 3'b100;
        rom_memory[17375] = 3'b110;
        rom_memory[17376] = 3'b110;
        rom_memory[17377] = 3'b110;
        rom_memory[17378] = 3'b110;
        rom_memory[17379] = 3'b110;
        rom_memory[17380] = 3'b110;
        rom_memory[17381] = 3'b110;
        rom_memory[17382] = 3'b111;
        rom_memory[17383] = 3'b110;
        rom_memory[17384] = 3'b100;
        rom_memory[17385] = 3'b110;
        rom_memory[17386] = 3'b110;
        rom_memory[17387] = 3'b110;
        rom_memory[17388] = 3'b110;
        rom_memory[17389] = 3'b110;
        rom_memory[17390] = 3'b111;
        rom_memory[17391] = 3'b111;
        rom_memory[17392] = 3'b111;
        rom_memory[17393] = 3'b110;
        rom_memory[17394] = 3'b110;
        rom_memory[17395] = 3'b110;
        rom_memory[17396] = 3'b110;
        rom_memory[17397] = 3'b110;
        rom_memory[17398] = 3'b110;
        rom_memory[17399] = 3'b110;
        rom_memory[17400] = 3'b110;
        rom_memory[17401] = 3'b110;
        rom_memory[17402] = 3'b110;
        rom_memory[17403] = 3'b110;
        rom_memory[17404] = 3'b110;
        rom_memory[17405] = 3'b110;
        rom_memory[17406] = 3'b110;
        rom_memory[17407] = 3'b111;
        rom_memory[17408] = 3'b111;
        rom_memory[17409] = 3'b111;
        rom_memory[17410] = 3'b111;
        rom_memory[17411] = 3'b111;
        rom_memory[17412] = 3'b110;
        rom_memory[17413] = 3'b110;
        rom_memory[17414] = 3'b110;
        rom_memory[17415] = 3'b110;
        rom_memory[17416] = 3'b111;
        rom_memory[17417] = 3'b111;
        rom_memory[17418] = 3'b111;
        rom_memory[17419] = 3'b111;
        rom_memory[17420] = 3'b111;
        rom_memory[17421] = 3'b111;
        rom_memory[17422] = 3'b111;
        rom_memory[17423] = 3'b111;
        rom_memory[17424] = 3'b111;
        rom_memory[17425] = 3'b111;
        rom_memory[17426] = 3'b111;
        rom_memory[17427] = 3'b111;
        rom_memory[17428] = 3'b111;
        rom_memory[17429] = 3'b111;
        rom_memory[17430] = 3'b111;
        rom_memory[17431] = 3'b111;
        rom_memory[17432] = 3'b111;
        rom_memory[17433] = 3'b111;
        rom_memory[17434] = 3'b111;
        rom_memory[17435] = 3'b111;
        rom_memory[17436] = 3'b111;
        rom_memory[17437] = 3'b111;
        rom_memory[17438] = 3'b111;
        rom_memory[17439] = 3'b111;
        rom_memory[17440] = 3'b111;
        rom_memory[17441] = 3'b111;
        rom_memory[17442] = 3'b111;
        rom_memory[17443] = 3'b111;
        rom_memory[17444] = 3'b111;
        rom_memory[17445] = 3'b111;
        rom_memory[17446] = 3'b111;
        rom_memory[17447] = 3'b111;
        rom_memory[17448] = 3'b111;
        rom_memory[17449] = 3'b111;
        rom_memory[17450] = 3'b111;
        rom_memory[17451] = 3'b111;
        rom_memory[17452] = 3'b111;
        rom_memory[17453] = 3'b111;
        rom_memory[17454] = 3'b111;
        rom_memory[17455] = 3'b111;
        rom_memory[17456] = 3'b111;
        rom_memory[17457] = 3'b111;
        rom_memory[17458] = 3'b111;
        rom_memory[17459] = 3'b111;
        rom_memory[17460] = 3'b111;
        rom_memory[17461] = 3'b111;
        rom_memory[17462] = 3'b111;
        rom_memory[17463] = 3'b110;
        rom_memory[17464] = 3'b111;
        rom_memory[17465] = 3'b110;
        rom_memory[17466] = 3'b110;
        rom_memory[17467] = 3'b110;
        rom_memory[17468] = 3'b111;
        rom_memory[17469] = 3'b111;
        rom_memory[17470] = 3'b110;
        rom_memory[17471] = 3'b110;
        rom_memory[17472] = 3'b110;
        rom_memory[17473] = 3'b110;
        rom_memory[17474] = 3'b110;
        rom_memory[17475] = 3'b110;
        rom_memory[17476] = 3'b110;
        rom_memory[17477] = 3'b110;
        rom_memory[17478] = 3'b110;
        rom_memory[17479] = 3'b110;
        rom_memory[17480] = 3'b110;
        rom_memory[17481] = 3'b110;
        rom_memory[17482] = 3'b110;
        rom_memory[17483] = 3'b110;
        rom_memory[17484] = 3'b110;
        rom_memory[17485] = 3'b110;
        rom_memory[17486] = 3'b110;
        rom_memory[17487] = 3'b110;
        rom_memory[17488] = 3'b110;
        rom_memory[17489] = 3'b110;
        rom_memory[17490] = 3'b110;
        rom_memory[17491] = 3'b110;
        rom_memory[17492] = 3'b110;
        rom_memory[17493] = 3'b110;
        rom_memory[17494] = 3'b110;
        rom_memory[17495] = 3'b110;
        rom_memory[17496] = 3'b110;
        rom_memory[17497] = 3'b110;
        rom_memory[17498] = 3'b110;
        rom_memory[17499] = 3'b110;
        rom_memory[17500] = 3'b110;
        rom_memory[17501] = 3'b110;
        rom_memory[17502] = 3'b110;
        rom_memory[17503] = 3'b110;
        rom_memory[17504] = 3'b110;
        rom_memory[17505] = 3'b110;
        rom_memory[17506] = 3'b110;
        rom_memory[17507] = 3'b110;
        rom_memory[17508] = 3'b110;
        rom_memory[17509] = 3'b110;
        rom_memory[17510] = 3'b110;
        rom_memory[17511] = 3'b110;
        rom_memory[17512] = 3'b110;
        rom_memory[17513] = 3'b110;
        rom_memory[17514] = 3'b110;
        rom_memory[17515] = 3'b110;
        rom_memory[17516] = 3'b110;
        rom_memory[17517] = 3'b110;
        rom_memory[17518] = 3'b110;
        rom_memory[17519] = 3'b110;
        rom_memory[17520] = 3'b110;
        rom_memory[17521] = 3'b110;
        rom_memory[17522] = 3'b110;
        rom_memory[17523] = 3'b110;
        rom_memory[17524] = 3'b110;
        rom_memory[17525] = 3'b110;
        rom_memory[17526] = 3'b110;
        rom_memory[17527] = 3'b110;
        rom_memory[17528] = 3'b110;
        rom_memory[17529] = 3'b110;
        rom_memory[17530] = 3'b110;
        rom_memory[17531] = 3'b110;
        rom_memory[17532] = 3'b110;
        rom_memory[17533] = 3'b110;
        rom_memory[17534] = 3'b110;
        rom_memory[17535] = 3'b110;
        rom_memory[17536] = 3'b110;
        rom_memory[17537] = 3'b110;
        rom_memory[17538] = 3'b110;
        rom_memory[17539] = 3'b110;
        rom_memory[17540] = 3'b110;
        rom_memory[17541] = 3'b110;
        rom_memory[17542] = 3'b110;
        rom_memory[17543] = 3'b110;
        rom_memory[17544] = 3'b110;
        rom_memory[17545] = 3'b110;
        rom_memory[17546] = 3'b110;
        rom_memory[17547] = 3'b110;
        rom_memory[17548] = 3'b110;
        rom_memory[17549] = 3'b110;
        rom_memory[17550] = 3'b110;
        rom_memory[17551] = 3'b110;
        rom_memory[17552] = 3'b110;
        rom_memory[17553] = 3'b110;
        rom_memory[17554] = 3'b111;
        rom_memory[17555] = 3'b111;
        rom_memory[17556] = 3'b111;
        rom_memory[17557] = 3'b111;
        rom_memory[17558] = 3'b111;
        rom_memory[17559] = 3'b111;
        rom_memory[17560] = 3'b111;
        rom_memory[17561] = 3'b111;
        rom_memory[17562] = 3'b111;
        rom_memory[17563] = 3'b111;
        rom_memory[17564] = 3'b111;
        rom_memory[17565] = 3'b110;
        rom_memory[17566] = 3'b100;
        rom_memory[17567] = 3'b100;
        rom_memory[17568] = 3'b100;
        rom_memory[17569] = 3'b100;
        rom_memory[17570] = 3'b100;
        rom_memory[17571] = 3'b100;
        rom_memory[17572] = 3'b100;
        rom_memory[17573] = 3'b100;
        rom_memory[17574] = 3'b100;
        rom_memory[17575] = 3'b100;
        rom_memory[17576] = 3'b100;
        rom_memory[17577] = 3'b100;
        rom_memory[17578] = 3'b100;
        rom_memory[17579] = 3'b100;
        rom_memory[17580] = 3'b100;
        rom_memory[17581] = 3'b100;
        rom_memory[17582] = 3'b100;
        rom_memory[17583] = 3'b100;
        rom_memory[17584] = 3'b110;
        rom_memory[17585] = 3'b110;
        rom_memory[17586] = 3'b110;
        rom_memory[17587] = 3'b110;
        rom_memory[17588] = 3'b100;
        rom_memory[17589] = 3'b110;
        rom_memory[17590] = 3'b110;
        rom_memory[17591] = 3'b100;
        rom_memory[17592] = 3'b110;
        rom_memory[17593] = 3'b110;
        rom_memory[17594] = 3'b110;
        rom_memory[17595] = 3'b110;
        rom_memory[17596] = 3'b110;
        rom_memory[17597] = 3'b110;
        rom_memory[17598] = 3'b110;
        rom_memory[17599] = 3'b110;
        rom_memory[17600] = 3'b110;
        rom_memory[17601] = 3'b110;
        rom_memory[17602] = 3'b110;
        rom_memory[17603] = 3'b110;
        rom_memory[17604] = 3'b110;
        rom_memory[17605] = 3'b110;
        rom_memory[17606] = 3'b110;
        rom_memory[17607] = 3'b110;
        rom_memory[17608] = 3'b110;
        rom_memory[17609] = 3'b110;
        rom_memory[17610] = 3'b000;
        rom_memory[17611] = 3'b000;
        rom_memory[17612] = 3'b000;
        rom_memory[17613] = 3'b000;
        rom_memory[17614] = 3'b000;
        rom_memory[17615] = 3'b100;
        rom_memory[17616] = 3'b110;
        rom_memory[17617] = 3'b110;
        rom_memory[17618] = 3'b110;
        rom_memory[17619] = 3'b110;
        rom_memory[17620] = 3'b110;
        rom_memory[17621] = 3'b110;
        rom_memory[17622] = 3'b110;
        rom_memory[17623] = 3'b110;
        rom_memory[17624] = 3'b110;
        rom_memory[17625] = 3'b110;
        rom_memory[17626] = 3'b110;
        rom_memory[17627] = 3'b110;
        rom_memory[17628] = 3'b110;
        rom_memory[17629] = 3'b100;
        rom_memory[17630] = 3'b110;
        rom_memory[17631] = 3'b111;
        rom_memory[17632] = 3'b111;
        rom_memory[17633] = 3'b111;
        rom_memory[17634] = 3'b111;
        rom_memory[17635] = 3'b110;
        rom_memory[17636] = 3'b110;
        rom_memory[17637] = 3'b110;
        rom_memory[17638] = 3'b110;
        rom_memory[17639] = 3'b110;
        rom_memory[17640] = 3'b110;
        rom_memory[17641] = 3'b110;
        rom_memory[17642] = 3'b110;
        rom_memory[17643] = 3'b110;
        rom_memory[17644] = 3'b110;
        rom_memory[17645] = 3'b110;
        rom_memory[17646] = 3'b110;
        rom_memory[17647] = 3'b111;
        rom_memory[17648] = 3'b110;
        rom_memory[17649] = 3'b110;
        rom_memory[17650] = 3'b110;
        rom_memory[17651] = 3'b110;
        rom_memory[17652] = 3'b111;
        rom_memory[17653] = 3'b111;
        rom_memory[17654] = 3'b111;
        rom_memory[17655] = 3'b110;
        rom_memory[17656] = 3'b110;
        rom_memory[17657] = 3'b111;
        rom_memory[17658] = 3'b111;
        rom_memory[17659] = 3'b111;
        rom_memory[17660] = 3'b111;
        rom_memory[17661] = 3'b111;
        rom_memory[17662] = 3'b111;
        rom_memory[17663] = 3'b111;
        rom_memory[17664] = 3'b111;
        rom_memory[17665] = 3'b111;
        rom_memory[17666] = 3'b111;
        rom_memory[17667] = 3'b111;
        rom_memory[17668] = 3'b111;
        rom_memory[17669] = 3'b111;
        rom_memory[17670] = 3'b111;
        rom_memory[17671] = 3'b111;
        rom_memory[17672] = 3'b111;
        rom_memory[17673] = 3'b111;
        rom_memory[17674] = 3'b111;
        rom_memory[17675] = 3'b111;
        rom_memory[17676] = 3'b111;
        rom_memory[17677] = 3'b111;
        rom_memory[17678] = 3'b111;
        rom_memory[17679] = 3'b111;
        rom_memory[17680] = 3'b111;
        rom_memory[17681] = 3'b111;
        rom_memory[17682] = 3'b111;
        rom_memory[17683] = 3'b111;
        rom_memory[17684] = 3'b111;
        rom_memory[17685] = 3'b111;
        rom_memory[17686] = 3'b111;
        rom_memory[17687] = 3'b111;
        rom_memory[17688] = 3'b111;
        rom_memory[17689] = 3'b111;
        rom_memory[17690] = 3'b111;
        rom_memory[17691] = 3'b111;
        rom_memory[17692] = 3'b111;
        rom_memory[17693] = 3'b111;
        rom_memory[17694] = 3'b111;
        rom_memory[17695] = 3'b111;
        rom_memory[17696] = 3'b111;
        rom_memory[17697] = 3'b111;
        rom_memory[17698] = 3'b111;
        rom_memory[17699] = 3'b111;
        rom_memory[17700] = 3'b111;
        rom_memory[17701] = 3'b111;
        rom_memory[17702] = 3'b111;
        rom_memory[17703] = 3'b111;
        rom_memory[17704] = 3'b111;
        rom_memory[17705] = 3'b111;
        rom_memory[17706] = 3'b110;
        rom_memory[17707] = 3'b110;
        rom_memory[17708] = 3'b111;
        rom_memory[17709] = 3'b111;
        rom_memory[17710] = 3'b110;
        rom_memory[17711] = 3'b110;
        rom_memory[17712] = 3'b110;
        rom_memory[17713] = 3'b110;
        rom_memory[17714] = 3'b110;
        rom_memory[17715] = 3'b110;
        rom_memory[17716] = 3'b110;
        rom_memory[17717] = 3'b110;
        rom_memory[17718] = 3'b110;
        rom_memory[17719] = 3'b110;
        rom_memory[17720] = 3'b110;
        rom_memory[17721] = 3'b110;
        rom_memory[17722] = 3'b110;
        rom_memory[17723] = 3'b110;
        rom_memory[17724] = 3'b110;
        rom_memory[17725] = 3'b110;
        rom_memory[17726] = 3'b110;
        rom_memory[17727] = 3'b110;
        rom_memory[17728] = 3'b110;
        rom_memory[17729] = 3'b110;
        rom_memory[17730] = 3'b110;
        rom_memory[17731] = 3'b110;
        rom_memory[17732] = 3'b110;
        rom_memory[17733] = 3'b110;
        rom_memory[17734] = 3'b110;
        rom_memory[17735] = 3'b110;
        rom_memory[17736] = 3'b110;
        rom_memory[17737] = 3'b110;
        rom_memory[17738] = 3'b110;
        rom_memory[17739] = 3'b110;
        rom_memory[17740] = 3'b110;
        rom_memory[17741] = 3'b110;
        rom_memory[17742] = 3'b110;
        rom_memory[17743] = 3'b110;
        rom_memory[17744] = 3'b110;
        rom_memory[17745] = 3'b110;
        rom_memory[17746] = 3'b110;
        rom_memory[17747] = 3'b110;
        rom_memory[17748] = 3'b110;
        rom_memory[17749] = 3'b110;
        rom_memory[17750] = 3'b110;
        rom_memory[17751] = 3'b110;
        rom_memory[17752] = 3'b110;
        rom_memory[17753] = 3'b110;
        rom_memory[17754] = 3'b110;
        rom_memory[17755] = 3'b110;
        rom_memory[17756] = 3'b110;
        rom_memory[17757] = 3'b110;
        rom_memory[17758] = 3'b110;
        rom_memory[17759] = 3'b110;
        rom_memory[17760] = 3'b110;
        rom_memory[17761] = 3'b110;
        rom_memory[17762] = 3'b110;
        rom_memory[17763] = 3'b110;
        rom_memory[17764] = 3'b110;
        rom_memory[17765] = 3'b110;
        rom_memory[17766] = 3'b110;
        rom_memory[17767] = 3'b110;
        rom_memory[17768] = 3'b110;
        rom_memory[17769] = 3'b110;
        rom_memory[17770] = 3'b110;
        rom_memory[17771] = 3'b110;
        rom_memory[17772] = 3'b110;
        rom_memory[17773] = 3'b110;
        rom_memory[17774] = 3'b110;
        rom_memory[17775] = 3'b110;
        rom_memory[17776] = 3'b110;
        rom_memory[17777] = 3'b110;
        rom_memory[17778] = 3'b110;
        rom_memory[17779] = 3'b110;
        rom_memory[17780] = 3'b110;
        rom_memory[17781] = 3'b110;
        rom_memory[17782] = 3'b110;
        rom_memory[17783] = 3'b110;
        rom_memory[17784] = 3'b110;
        rom_memory[17785] = 3'b110;
        rom_memory[17786] = 3'b110;
        rom_memory[17787] = 3'b110;
        rom_memory[17788] = 3'b110;
        rom_memory[17789] = 3'b110;
        rom_memory[17790] = 3'b110;
        rom_memory[17791] = 3'b110;
        rom_memory[17792] = 3'b110;
        rom_memory[17793] = 3'b111;
        rom_memory[17794] = 3'b111;
        rom_memory[17795] = 3'b111;
        rom_memory[17796] = 3'b111;
        rom_memory[17797] = 3'b111;
        rom_memory[17798] = 3'b111;
        rom_memory[17799] = 3'b111;
        rom_memory[17800] = 3'b111;
        rom_memory[17801] = 3'b111;
        rom_memory[17802] = 3'b111;
        rom_memory[17803] = 3'b111;
        rom_memory[17804] = 3'b111;
        rom_memory[17805] = 3'b100;
        rom_memory[17806] = 3'b100;
        rom_memory[17807] = 3'b100;
        rom_memory[17808] = 3'b100;
        rom_memory[17809] = 3'b100;
        rom_memory[17810] = 3'b100;
        rom_memory[17811] = 3'b100;
        rom_memory[17812] = 3'b110;
        rom_memory[17813] = 3'b110;
        rom_memory[17814] = 3'b110;
        rom_memory[17815] = 3'b100;
        rom_memory[17816] = 3'b100;
        rom_memory[17817] = 3'b100;
        rom_memory[17818] = 3'b100;
        rom_memory[17819] = 3'b100;
        rom_memory[17820] = 3'b100;
        rom_memory[17821] = 3'b100;
        rom_memory[17822] = 3'b100;
        rom_memory[17823] = 3'b100;
        rom_memory[17824] = 3'b100;
        rom_memory[17825] = 3'b110;
        rom_memory[17826] = 3'b110;
        rom_memory[17827] = 3'b100;
        rom_memory[17828] = 3'b100;
        rom_memory[17829] = 3'b110;
        rom_memory[17830] = 3'b110;
        rom_memory[17831] = 3'b110;
        rom_memory[17832] = 3'b110;
        rom_memory[17833] = 3'b110;
        rom_memory[17834] = 3'b110;
        rom_memory[17835] = 3'b110;
        rom_memory[17836] = 3'b110;
        rom_memory[17837] = 3'b110;
        rom_memory[17838] = 3'b110;
        rom_memory[17839] = 3'b110;
        rom_memory[17840] = 3'b110;
        rom_memory[17841] = 3'b110;
        rom_memory[17842] = 3'b110;
        rom_memory[17843] = 3'b110;
        rom_memory[17844] = 3'b110;
        rom_memory[17845] = 3'b110;
        rom_memory[17846] = 3'b110;
        rom_memory[17847] = 3'b110;
        rom_memory[17848] = 3'b110;
        rom_memory[17849] = 3'b110;
        rom_memory[17850] = 3'b110;
        rom_memory[17851] = 3'b000;
        rom_memory[17852] = 3'b000;
        rom_memory[17853] = 3'b000;
        rom_memory[17854] = 3'b000;
        rom_memory[17855] = 3'b000;
        rom_memory[17856] = 3'b100;
        rom_memory[17857] = 3'b110;
        rom_memory[17858] = 3'b110;
        rom_memory[17859] = 3'b110;
        rom_memory[17860] = 3'b110;
        rom_memory[17861] = 3'b110;
        rom_memory[17862] = 3'b110;
        rom_memory[17863] = 3'b110;
        rom_memory[17864] = 3'b110;
        rom_memory[17865] = 3'b110;
        rom_memory[17866] = 3'b110;
        rom_memory[17867] = 3'b110;
        rom_memory[17868] = 3'b110;
        rom_memory[17869] = 3'b110;
        rom_memory[17870] = 3'b100;
        rom_memory[17871] = 3'b110;
        rom_memory[17872] = 3'b111;
        rom_memory[17873] = 3'b111;
        rom_memory[17874] = 3'b111;
        rom_memory[17875] = 3'b110;
        rom_memory[17876] = 3'b110;
        rom_memory[17877] = 3'b110;
        rom_memory[17878] = 3'b110;
        rom_memory[17879] = 3'b110;
        rom_memory[17880] = 3'b110;
        rom_memory[17881] = 3'b110;
        rom_memory[17882] = 3'b110;
        rom_memory[17883] = 3'b110;
        rom_memory[17884] = 3'b110;
        rom_memory[17885] = 3'b110;
        rom_memory[17886] = 3'b110;
        rom_memory[17887] = 3'b110;
        rom_memory[17888] = 3'b110;
        rom_memory[17889] = 3'b110;
        rom_memory[17890] = 3'b111;
        rom_memory[17891] = 3'b111;
        rom_memory[17892] = 3'b111;
        rom_memory[17893] = 3'b111;
        rom_memory[17894] = 3'b111;
        rom_memory[17895] = 3'b110;
        rom_memory[17896] = 3'b110;
        rom_memory[17897] = 3'b111;
        rom_memory[17898] = 3'b111;
        rom_memory[17899] = 3'b111;
        rom_memory[17900] = 3'b111;
        rom_memory[17901] = 3'b111;
        rom_memory[17902] = 3'b111;
        rom_memory[17903] = 3'b111;
        rom_memory[17904] = 3'b111;
        rom_memory[17905] = 3'b111;
        rom_memory[17906] = 3'b111;
        rom_memory[17907] = 3'b111;
        rom_memory[17908] = 3'b111;
        rom_memory[17909] = 3'b111;
        rom_memory[17910] = 3'b111;
        rom_memory[17911] = 3'b111;
        rom_memory[17912] = 3'b111;
        rom_memory[17913] = 3'b111;
        rom_memory[17914] = 3'b111;
        rom_memory[17915] = 3'b111;
        rom_memory[17916] = 3'b111;
        rom_memory[17917] = 3'b111;
        rom_memory[17918] = 3'b111;
        rom_memory[17919] = 3'b111;
        rom_memory[17920] = 3'b111;
        rom_memory[17921] = 3'b111;
        rom_memory[17922] = 3'b111;
        rom_memory[17923] = 3'b111;
        rom_memory[17924] = 3'b111;
        rom_memory[17925] = 3'b111;
        rom_memory[17926] = 3'b111;
        rom_memory[17927] = 3'b111;
        rom_memory[17928] = 3'b111;
        rom_memory[17929] = 3'b111;
        rom_memory[17930] = 3'b111;
        rom_memory[17931] = 3'b111;
        rom_memory[17932] = 3'b111;
        rom_memory[17933] = 3'b111;
        rom_memory[17934] = 3'b111;
        rom_memory[17935] = 3'b111;
        rom_memory[17936] = 3'b111;
        rom_memory[17937] = 3'b111;
        rom_memory[17938] = 3'b111;
        rom_memory[17939] = 3'b111;
        rom_memory[17940] = 3'b111;
        rom_memory[17941] = 3'b111;
        rom_memory[17942] = 3'b111;
        rom_memory[17943] = 3'b111;
        rom_memory[17944] = 3'b111;
        rom_memory[17945] = 3'b111;
        rom_memory[17946] = 3'b110;
        rom_memory[17947] = 3'b110;
        rom_memory[17948] = 3'b110;
        rom_memory[17949] = 3'b111;
        rom_memory[17950] = 3'b110;
        rom_memory[17951] = 3'b110;
        rom_memory[17952] = 3'b110;
        rom_memory[17953] = 3'b110;
        rom_memory[17954] = 3'b110;
        rom_memory[17955] = 3'b110;
        rom_memory[17956] = 3'b110;
        rom_memory[17957] = 3'b110;
        rom_memory[17958] = 3'b110;
        rom_memory[17959] = 3'b110;
        rom_memory[17960] = 3'b110;
        rom_memory[17961] = 3'b110;
        rom_memory[17962] = 3'b110;
        rom_memory[17963] = 3'b110;
        rom_memory[17964] = 3'b110;
        rom_memory[17965] = 3'b110;
        rom_memory[17966] = 3'b110;
        rom_memory[17967] = 3'b110;
        rom_memory[17968] = 3'b110;
        rom_memory[17969] = 3'b110;
        rom_memory[17970] = 3'b110;
        rom_memory[17971] = 3'b110;
        rom_memory[17972] = 3'b110;
        rom_memory[17973] = 3'b110;
        rom_memory[17974] = 3'b110;
        rom_memory[17975] = 3'b110;
        rom_memory[17976] = 3'b110;
        rom_memory[17977] = 3'b110;
        rom_memory[17978] = 3'b110;
        rom_memory[17979] = 3'b110;
        rom_memory[17980] = 3'b110;
        rom_memory[17981] = 3'b110;
        rom_memory[17982] = 3'b110;
        rom_memory[17983] = 3'b110;
        rom_memory[17984] = 3'b110;
        rom_memory[17985] = 3'b110;
        rom_memory[17986] = 3'b110;
        rom_memory[17987] = 3'b110;
        rom_memory[17988] = 3'b110;
        rom_memory[17989] = 3'b110;
        rom_memory[17990] = 3'b110;
        rom_memory[17991] = 3'b110;
        rom_memory[17992] = 3'b110;
        rom_memory[17993] = 3'b110;
        rom_memory[17994] = 3'b110;
        rom_memory[17995] = 3'b110;
        rom_memory[17996] = 3'b110;
        rom_memory[17997] = 3'b110;
        rom_memory[17998] = 3'b110;
        rom_memory[17999] = 3'b110;
        rom_memory[18000] = 3'b110;
        rom_memory[18001] = 3'b110;
        rom_memory[18002] = 3'b110;
        rom_memory[18003] = 3'b110;
        rom_memory[18004] = 3'b110;
        rom_memory[18005] = 3'b110;
        rom_memory[18006] = 3'b110;
        rom_memory[18007] = 3'b110;
        rom_memory[18008] = 3'b110;
        rom_memory[18009] = 3'b110;
        rom_memory[18010] = 3'b110;
        rom_memory[18011] = 3'b110;
        rom_memory[18012] = 3'b110;
        rom_memory[18013] = 3'b110;
        rom_memory[18014] = 3'b110;
        rom_memory[18015] = 3'b110;
        rom_memory[18016] = 3'b110;
        rom_memory[18017] = 3'b110;
        rom_memory[18018] = 3'b110;
        rom_memory[18019] = 3'b110;
        rom_memory[18020] = 3'b110;
        rom_memory[18021] = 3'b110;
        rom_memory[18022] = 3'b110;
        rom_memory[18023] = 3'b110;
        rom_memory[18024] = 3'b110;
        rom_memory[18025] = 3'b110;
        rom_memory[18026] = 3'b110;
        rom_memory[18027] = 3'b110;
        rom_memory[18028] = 3'b110;
        rom_memory[18029] = 3'b110;
        rom_memory[18030] = 3'b110;
        rom_memory[18031] = 3'b111;
        rom_memory[18032] = 3'b111;
        rom_memory[18033] = 3'b111;
        rom_memory[18034] = 3'b111;
        rom_memory[18035] = 3'b111;
        rom_memory[18036] = 3'b111;
        rom_memory[18037] = 3'b111;
        rom_memory[18038] = 3'b111;
        rom_memory[18039] = 3'b111;
        rom_memory[18040] = 3'b111;
        rom_memory[18041] = 3'b111;
        rom_memory[18042] = 3'b111;
        rom_memory[18043] = 3'b111;
        rom_memory[18044] = 3'b111;
        rom_memory[18045] = 3'b100;
        rom_memory[18046] = 3'b100;
        rom_memory[18047] = 3'b100;
        rom_memory[18048] = 3'b100;
        rom_memory[18049] = 3'b100;
        rom_memory[18050] = 3'b100;
        rom_memory[18051] = 3'b100;
        rom_memory[18052] = 3'b110;
        rom_memory[18053] = 3'b110;
        rom_memory[18054] = 3'b110;
        rom_memory[18055] = 3'b100;
        rom_memory[18056] = 3'b100;
        rom_memory[18057] = 3'b110;
        rom_memory[18058] = 3'b110;
        rom_memory[18059] = 3'b110;
        rom_memory[18060] = 3'b100;
        rom_memory[18061] = 3'b110;
        rom_memory[18062] = 3'b110;
        rom_memory[18063] = 3'b110;
        rom_memory[18064] = 3'b110;
        rom_memory[18065] = 3'b110;
        rom_memory[18066] = 3'b110;
        rom_memory[18067] = 3'b110;
        rom_memory[18068] = 3'b110;
        rom_memory[18069] = 3'b110;
        rom_memory[18070] = 3'b100;
        rom_memory[18071] = 3'b100;
        rom_memory[18072] = 3'b110;
        rom_memory[18073] = 3'b110;
        rom_memory[18074] = 3'b110;
        rom_memory[18075] = 3'b110;
        rom_memory[18076] = 3'b110;
        rom_memory[18077] = 3'b110;
        rom_memory[18078] = 3'b110;
        rom_memory[18079] = 3'b110;
        rom_memory[18080] = 3'b110;
        rom_memory[18081] = 3'b110;
        rom_memory[18082] = 3'b110;
        rom_memory[18083] = 3'b110;
        rom_memory[18084] = 3'b110;
        rom_memory[18085] = 3'b110;
        rom_memory[18086] = 3'b110;
        rom_memory[18087] = 3'b110;
        rom_memory[18088] = 3'b110;
        rom_memory[18089] = 3'b110;
        rom_memory[18090] = 3'b110;
        rom_memory[18091] = 3'b110;
        rom_memory[18092] = 3'b000;
        rom_memory[18093] = 3'b000;
        rom_memory[18094] = 3'b100;
        rom_memory[18095] = 3'b000;
        rom_memory[18096] = 3'b000;
        rom_memory[18097] = 3'b100;
        rom_memory[18098] = 3'b110;
        rom_memory[18099] = 3'b110;
        rom_memory[18100] = 3'b110;
        rom_memory[18101] = 3'b110;
        rom_memory[18102] = 3'b110;
        rom_memory[18103] = 3'b110;
        rom_memory[18104] = 3'b110;
        rom_memory[18105] = 3'b110;
        rom_memory[18106] = 3'b110;
        rom_memory[18107] = 3'b110;
        rom_memory[18108] = 3'b110;
        rom_memory[18109] = 3'b110;
        rom_memory[18110] = 3'b110;
        rom_memory[18111] = 3'b000;
        rom_memory[18112] = 3'b110;
        rom_memory[18113] = 3'b111;
        rom_memory[18114] = 3'b111;
        rom_memory[18115] = 3'b111;
        rom_memory[18116] = 3'b110;
        rom_memory[18117] = 3'b110;
        rom_memory[18118] = 3'b110;
        rom_memory[18119] = 3'b110;
        rom_memory[18120] = 3'b110;
        rom_memory[18121] = 3'b110;
        rom_memory[18122] = 3'b110;
        rom_memory[18123] = 3'b110;
        rom_memory[18124] = 3'b110;
        rom_memory[18125] = 3'b110;
        rom_memory[18126] = 3'b110;
        rom_memory[18127] = 3'b110;
        rom_memory[18128] = 3'b110;
        rom_memory[18129] = 3'b110;
        rom_memory[18130] = 3'b110;
        rom_memory[18131] = 3'b111;
        rom_memory[18132] = 3'b111;
        rom_memory[18133] = 3'b111;
        rom_memory[18134] = 3'b110;
        rom_memory[18135] = 3'b110;
        rom_memory[18136] = 3'b110;
        rom_memory[18137] = 3'b110;
        rom_memory[18138] = 3'b111;
        rom_memory[18139] = 3'b111;
        rom_memory[18140] = 3'b111;
        rom_memory[18141] = 3'b111;
        rom_memory[18142] = 3'b111;
        rom_memory[18143] = 3'b111;
        rom_memory[18144] = 3'b111;
        rom_memory[18145] = 3'b111;
        rom_memory[18146] = 3'b111;
        rom_memory[18147] = 3'b111;
        rom_memory[18148] = 3'b111;
        rom_memory[18149] = 3'b111;
        rom_memory[18150] = 3'b111;
        rom_memory[18151] = 3'b111;
        rom_memory[18152] = 3'b111;
        rom_memory[18153] = 3'b111;
        rom_memory[18154] = 3'b111;
        rom_memory[18155] = 3'b111;
        rom_memory[18156] = 3'b111;
        rom_memory[18157] = 3'b111;
        rom_memory[18158] = 3'b111;
        rom_memory[18159] = 3'b111;
        rom_memory[18160] = 3'b111;
        rom_memory[18161] = 3'b111;
        rom_memory[18162] = 3'b111;
        rom_memory[18163] = 3'b111;
        rom_memory[18164] = 3'b111;
        rom_memory[18165] = 3'b111;
        rom_memory[18166] = 3'b111;
        rom_memory[18167] = 3'b111;
        rom_memory[18168] = 3'b111;
        rom_memory[18169] = 3'b111;
        rom_memory[18170] = 3'b111;
        rom_memory[18171] = 3'b111;
        rom_memory[18172] = 3'b111;
        rom_memory[18173] = 3'b111;
        rom_memory[18174] = 3'b111;
        rom_memory[18175] = 3'b111;
        rom_memory[18176] = 3'b111;
        rom_memory[18177] = 3'b111;
        rom_memory[18178] = 3'b111;
        rom_memory[18179] = 3'b111;
        rom_memory[18180] = 3'b111;
        rom_memory[18181] = 3'b111;
        rom_memory[18182] = 3'b111;
        rom_memory[18183] = 3'b111;
        rom_memory[18184] = 3'b111;
        rom_memory[18185] = 3'b111;
        rom_memory[18186] = 3'b111;
        rom_memory[18187] = 3'b110;
        rom_memory[18188] = 3'b110;
        rom_memory[18189] = 3'b111;
        rom_memory[18190] = 3'b111;
        rom_memory[18191] = 3'b110;
        rom_memory[18192] = 3'b110;
        rom_memory[18193] = 3'b110;
        rom_memory[18194] = 3'b110;
        rom_memory[18195] = 3'b110;
        rom_memory[18196] = 3'b110;
        rom_memory[18197] = 3'b110;
        rom_memory[18198] = 3'b110;
        rom_memory[18199] = 3'b110;
        rom_memory[18200] = 3'b110;
        rom_memory[18201] = 3'b110;
        rom_memory[18202] = 3'b110;
        rom_memory[18203] = 3'b110;
        rom_memory[18204] = 3'b110;
        rom_memory[18205] = 3'b110;
        rom_memory[18206] = 3'b110;
        rom_memory[18207] = 3'b110;
        rom_memory[18208] = 3'b110;
        rom_memory[18209] = 3'b110;
        rom_memory[18210] = 3'b110;
        rom_memory[18211] = 3'b110;
        rom_memory[18212] = 3'b110;
        rom_memory[18213] = 3'b110;
        rom_memory[18214] = 3'b110;
        rom_memory[18215] = 3'b110;
        rom_memory[18216] = 3'b110;
        rom_memory[18217] = 3'b110;
        rom_memory[18218] = 3'b110;
        rom_memory[18219] = 3'b110;
        rom_memory[18220] = 3'b110;
        rom_memory[18221] = 3'b110;
        rom_memory[18222] = 3'b110;
        rom_memory[18223] = 3'b110;
        rom_memory[18224] = 3'b110;
        rom_memory[18225] = 3'b110;
        rom_memory[18226] = 3'b110;
        rom_memory[18227] = 3'b110;
        rom_memory[18228] = 3'b110;
        rom_memory[18229] = 3'b110;
        rom_memory[18230] = 3'b110;
        rom_memory[18231] = 3'b110;
        rom_memory[18232] = 3'b110;
        rom_memory[18233] = 3'b110;
        rom_memory[18234] = 3'b110;
        rom_memory[18235] = 3'b110;
        rom_memory[18236] = 3'b110;
        rom_memory[18237] = 3'b110;
        rom_memory[18238] = 3'b110;
        rom_memory[18239] = 3'b110;
        rom_memory[18240] = 3'b110;
        rom_memory[18241] = 3'b110;
        rom_memory[18242] = 3'b110;
        rom_memory[18243] = 3'b110;
        rom_memory[18244] = 3'b110;
        rom_memory[18245] = 3'b110;
        rom_memory[18246] = 3'b110;
        rom_memory[18247] = 3'b110;
        rom_memory[18248] = 3'b110;
        rom_memory[18249] = 3'b110;
        rom_memory[18250] = 3'b110;
        rom_memory[18251] = 3'b110;
        rom_memory[18252] = 3'b110;
        rom_memory[18253] = 3'b110;
        rom_memory[18254] = 3'b110;
        rom_memory[18255] = 3'b110;
        rom_memory[18256] = 3'b110;
        rom_memory[18257] = 3'b110;
        rom_memory[18258] = 3'b110;
        rom_memory[18259] = 3'b110;
        rom_memory[18260] = 3'b110;
        rom_memory[18261] = 3'b110;
        rom_memory[18262] = 3'b110;
        rom_memory[18263] = 3'b110;
        rom_memory[18264] = 3'b110;
        rom_memory[18265] = 3'b110;
        rom_memory[18266] = 3'b110;
        rom_memory[18267] = 3'b110;
        rom_memory[18268] = 3'b110;
        rom_memory[18269] = 3'b110;
        rom_memory[18270] = 3'b110;
        rom_memory[18271] = 3'b111;
        rom_memory[18272] = 3'b111;
        rom_memory[18273] = 3'b111;
        rom_memory[18274] = 3'b111;
        rom_memory[18275] = 3'b111;
        rom_memory[18276] = 3'b111;
        rom_memory[18277] = 3'b111;
        rom_memory[18278] = 3'b111;
        rom_memory[18279] = 3'b111;
        rom_memory[18280] = 3'b111;
        rom_memory[18281] = 3'b111;
        rom_memory[18282] = 3'b111;
        rom_memory[18283] = 3'b111;
        rom_memory[18284] = 3'b111;
        rom_memory[18285] = 3'b100;
        rom_memory[18286] = 3'b100;
        rom_memory[18287] = 3'b100;
        rom_memory[18288] = 3'b100;
        rom_memory[18289] = 3'b100;
        rom_memory[18290] = 3'b100;
        rom_memory[18291] = 3'b110;
        rom_memory[18292] = 3'b110;
        rom_memory[18293] = 3'b110;
        rom_memory[18294] = 3'b100;
        rom_memory[18295] = 3'b100;
        rom_memory[18296] = 3'b110;
        rom_memory[18297] = 3'b110;
        rom_memory[18298] = 3'b110;
        rom_memory[18299] = 3'b110;
        rom_memory[18300] = 3'b100;
        rom_memory[18301] = 3'b110;
        rom_memory[18302] = 3'b110;
        rom_memory[18303] = 3'b110;
        rom_memory[18304] = 3'b110;
        rom_memory[18305] = 3'b110;
        rom_memory[18306] = 3'b100;
        rom_memory[18307] = 3'b110;
        rom_memory[18308] = 3'b110;
        rom_memory[18309] = 3'b110;
        rom_memory[18310] = 3'b110;
        rom_memory[18311] = 3'b110;
        rom_memory[18312] = 3'b110;
        rom_memory[18313] = 3'b110;
        rom_memory[18314] = 3'b110;
        rom_memory[18315] = 3'b110;
        rom_memory[18316] = 3'b110;
        rom_memory[18317] = 3'b110;
        rom_memory[18318] = 3'b110;
        rom_memory[18319] = 3'b110;
        rom_memory[18320] = 3'b110;
        rom_memory[18321] = 3'b110;
        rom_memory[18322] = 3'b100;
        rom_memory[18323] = 3'b110;
        rom_memory[18324] = 3'b110;
        rom_memory[18325] = 3'b110;
        rom_memory[18326] = 3'b110;
        rom_memory[18327] = 3'b110;
        rom_memory[18328] = 3'b110;
        rom_memory[18329] = 3'b110;
        rom_memory[18330] = 3'b110;
        rom_memory[18331] = 3'b110;
        rom_memory[18332] = 3'b110;
        rom_memory[18333] = 3'b000;
        rom_memory[18334] = 3'b000;
        rom_memory[18335] = 3'b110;
        rom_memory[18336] = 3'b000;
        rom_memory[18337] = 3'b000;
        rom_memory[18338] = 3'b100;
        rom_memory[18339] = 3'b110;
        rom_memory[18340] = 3'b100;
        rom_memory[18341] = 3'b110;
        rom_memory[18342] = 3'b110;
        rom_memory[18343] = 3'b110;
        rom_memory[18344] = 3'b100;
        rom_memory[18345] = 3'b110;
        rom_memory[18346] = 3'b110;
        rom_memory[18347] = 3'b100;
        rom_memory[18348] = 3'b100;
        rom_memory[18349] = 3'b110;
        rom_memory[18350] = 3'b110;
        rom_memory[18351] = 3'b110;
        rom_memory[18352] = 3'b100;
        rom_memory[18353] = 3'b111;
        rom_memory[18354] = 3'b111;
        rom_memory[18355] = 3'b111;
        rom_memory[18356] = 3'b111;
        rom_memory[18357] = 3'b110;
        rom_memory[18358] = 3'b110;
        rom_memory[18359] = 3'b110;
        rom_memory[18360] = 3'b110;
        rom_memory[18361] = 3'b110;
        rom_memory[18362] = 3'b110;
        rom_memory[18363] = 3'b110;
        rom_memory[18364] = 3'b110;
        rom_memory[18365] = 3'b110;
        rom_memory[18366] = 3'b110;
        rom_memory[18367] = 3'b110;
        rom_memory[18368] = 3'b111;
        rom_memory[18369] = 3'b110;
        rom_memory[18370] = 3'b110;
        rom_memory[18371] = 3'b110;
        rom_memory[18372] = 3'b110;
        rom_memory[18373] = 3'b111;
        rom_memory[18374] = 3'b110;
        rom_memory[18375] = 3'b111;
        rom_memory[18376] = 3'b110;
        rom_memory[18377] = 3'b110;
        rom_memory[18378] = 3'b110;
        rom_memory[18379] = 3'b110;
        rom_memory[18380] = 3'b111;
        rom_memory[18381] = 3'b111;
        rom_memory[18382] = 3'b111;
        rom_memory[18383] = 3'b111;
        rom_memory[18384] = 3'b111;
        rom_memory[18385] = 3'b111;
        rom_memory[18386] = 3'b111;
        rom_memory[18387] = 3'b111;
        rom_memory[18388] = 3'b111;
        rom_memory[18389] = 3'b111;
        rom_memory[18390] = 3'b111;
        rom_memory[18391] = 3'b111;
        rom_memory[18392] = 3'b111;
        rom_memory[18393] = 3'b111;
        rom_memory[18394] = 3'b111;
        rom_memory[18395] = 3'b111;
        rom_memory[18396] = 3'b111;
        rom_memory[18397] = 3'b111;
        rom_memory[18398] = 3'b111;
        rom_memory[18399] = 3'b111;
        rom_memory[18400] = 3'b111;
        rom_memory[18401] = 3'b111;
        rom_memory[18402] = 3'b111;
        rom_memory[18403] = 3'b111;
        rom_memory[18404] = 3'b111;
        rom_memory[18405] = 3'b111;
        rom_memory[18406] = 3'b111;
        rom_memory[18407] = 3'b111;
        rom_memory[18408] = 3'b111;
        rom_memory[18409] = 3'b111;
        rom_memory[18410] = 3'b111;
        rom_memory[18411] = 3'b111;
        rom_memory[18412] = 3'b111;
        rom_memory[18413] = 3'b111;
        rom_memory[18414] = 3'b111;
        rom_memory[18415] = 3'b111;
        rom_memory[18416] = 3'b111;
        rom_memory[18417] = 3'b111;
        rom_memory[18418] = 3'b111;
        rom_memory[18419] = 3'b111;
        rom_memory[18420] = 3'b111;
        rom_memory[18421] = 3'b111;
        rom_memory[18422] = 3'b111;
        rom_memory[18423] = 3'b111;
        rom_memory[18424] = 3'b111;
        rom_memory[18425] = 3'b111;
        rom_memory[18426] = 3'b111;
        rom_memory[18427] = 3'b110;
        rom_memory[18428] = 3'b110;
        rom_memory[18429] = 3'b111;
        rom_memory[18430] = 3'b111;
        rom_memory[18431] = 3'b110;
        rom_memory[18432] = 3'b110;
        rom_memory[18433] = 3'b110;
        rom_memory[18434] = 3'b110;
        rom_memory[18435] = 3'b110;
        rom_memory[18436] = 3'b110;
        rom_memory[18437] = 3'b110;
        rom_memory[18438] = 3'b110;
        rom_memory[18439] = 3'b110;
        rom_memory[18440] = 3'b110;
        rom_memory[18441] = 3'b110;
        rom_memory[18442] = 3'b110;
        rom_memory[18443] = 3'b110;
        rom_memory[18444] = 3'b110;
        rom_memory[18445] = 3'b110;
        rom_memory[18446] = 3'b110;
        rom_memory[18447] = 3'b110;
        rom_memory[18448] = 3'b110;
        rom_memory[18449] = 3'b110;
        rom_memory[18450] = 3'b110;
        rom_memory[18451] = 3'b110;
        rom_memory[18452] = 3'b110;
        rom_memory[18453] = 3'b110;
        rom_memory[18454] = 3'b110;
        rom_memory[18455] = 3'b110;
        rom_memory[18456] = 3'b110;
        rom_memory[18457] = 3'b110;
        rom_memory[18458] = 3'b110;
        rom_memory[18459] = 3'b110;
        rom_memory[18460] = 3'b110;
        rom_memory[18461] = 3'b110;
        rom_memory[18462] = 3'b110;
        rom_memory[18463] = 3'b110;
        rom_memory[18464] = 3'b110;
        rom_memory[18465] = 3'b110;
        rom_memory[18466] = 3'b110;
        rom_memory[18467] = 3'b110;
        rom_memory[18468] = 3'b110;
        rom_memory[18469] = 3'b110;
        rom_memory[18470] = 3'b110;
        rom_memory[18471] = 3'b110;
        rom_memory[18472] = 3'b110;
        rom_memory[18473] = 3'b110;
        rom_memory[18474] = 3'b110;
        rom_memory[18475] = 3'b110;
        rom_memory[18476] = 3'b110;
        rom_memory[18477] = 3'b110;
        rom_memory[18478] = 3'b110;
        rom_memory[18479] = 3'b110;
        rom_memory[18480] = 3'b110;
        rom_memory[18481] = 3'b110;
        rom_memory[18482] = 3'b110;
        rom_memory[18483] = 3'b110;
        rom_memory[18484] = 3'b110;
        rom_memory[18485] = 3'b110;
        rom_memory[18486] = 3'b110;
        rom_memory[18487] = 3'b110;
        rom_memory[18488] = 3'b110;
        rom_memory[18489] = 3'b110;
        rom_memory[18490] = 3'b110;
        rom_memory[18491] = 3'b110;
        rom_memory[18492] = 3'b110;
        rom_memory[18493] = 3'b110;
        rom_memory[18494] = 3'b110;
        rom_memory[18495] = 3'b110;
        rom_memory[18496] = 3'b110;
        rom_memory[18497] = 3'b110;
        rom_memory[18498] = 3'b110;
        rom_memory[18499] = 3'b110;
        rom_memory[18500] = 3'b110;
        rom_memory[18501] = 3'b110;
        rom_memory[18502] = 3'b110;
        rom_memory[18503] = 3'b110;
        rom_memory[18504] = 3'b110;
        rom_memory[18505] = 3'b110;
        rom_memory[18506] = 3'b110;
        rom_memory[18507] = 3'b110;
        rom_memory[18508] = 3'b110;
        rom_memory[18509] = 3'b110;
        rom_memory[18510] = 3'b111;
        rom_memory[18511] = 3'b111;
        rom_memory[18512] = 3'b111;
        rom_memory[18513] = 3'b111;
        rom_memory[18514] = 3'b111;
        rom_memory[18515] = 3'b111;
        rom_memory[18516] = 3'b111;
        rom_memory[18517] = 3'b111;
        rom_memory[18518] = 3'b111;
        rom_memory[18519] = 3'b111;
        rom_memory[18520] = 3'b111;
        rom_memory[18521] = 3'b111;
        rom_memory[18522] = 3'b111;
        rom_memory[18523] = 3'b111;
        rom_memory[18524] = 3'b111;
        rom_memory[18525] = 3'b110;
        rom_memory[18526] = 3'b100;
        rom_memory[18527] = 3'b100;
        rom_memory[18528] = 3'b100;
        rom_memory[18529] = 3'b100;
        rom_memory[18530] = 3'b100;
        rom_memory[18531] = 3'b100;
        rom_memory[18532] = 3'b110;
        rom_memory[18533] = 3'b100;
        rom_memory[18534] = 3'b100;
        rom_memory[18535] = 3'b110;
        rom_memory[18536] = 3'b100;
        rom_memory[18537] = 3'b110;
        rom_memory[18538] = 3'b110;
        rom_memory[18539] = 3'b110;
        rom_memory[18540] = 3'b100;
        rom_memory[18541] = 3'b100;
        rom_memory[18542] = 3'b100;
        rom_memory[18543] = 3'b100;
        rom_memory[18544] = 3'b110;
        rom_memory[18545] = 3'b110;
        rom_memory[18546] = 3'b110;
        rom_memory[18547] = 3'b110;
        rom_memory[18548] = 3'b110;
        rom_memory[18549] = 3'b110;
        rom_memory[18550] = 3'b110;
        rom_memory[18551] = 3'b110;
        rom_memory[18552] = 3'b110;
        rom_memory[18553] = 3'b110;
        rom_memory[18554] = 3'b110;
        rom_memory[18555] = 3'b110;
        rom_memory[18556] = 3'b110;
        rom_memory[18557] = 3'b110;
        rom_memory[18558] = 3'b110;
        rom_memory[18559] = 3'b110;
        rom_memory[18560] = 3'b110;
        rom_memory[18561] = 3'b110;
        rom_memory[18562] = 3'b110;
        rom_memory[18563] = 3'b110;
        rom_memory[18564] = 3'b110;
        rom_memory[18565] = 3'b110;
        rom_memory[18566] = 3'b110;
        rom_memory[18567] = 3'b110;
        rom_memory[18568] = 3'b110;
        rom_memory[18569] = 3'b110;
        rom_memory[18570] = 3'b110;
        rom_memory[18571] = 3'b110;
        rom_memory[18572] = 3'b110;
        rom_memory[18573] = 3'b110;
        rom_memory[18574] = 3'b000;
        rom_memory[18575] = 3'b000;
        rom_memory[18576] = 3'b100;
        rom_memory[18577] = 3'b000;
        rom_memory[18578] = 3'b000;
        rom_memory[18579] = 3'b100;
        rom_memory[18580] = 3'b100;
        rom_memory[18581] = 3'b100;
        rom_memory[18582] = 3'b110;
        rom_memory[18583] = 3'b110;
        rom_memory[18584] = 3'b110;
        rom_memory[18585] = 3'b000;
        rom_memory[18586] = 3'b100;
        rom_memory[18587] = 3'b110;
        rom_memory[18588] = 3'b100;
        rom_memory[18589] = 3'b100;
        rom_memory[18590] = 3'b110;
        rom_memory[18591] = 3'b111;
        rom_memory[18592] = 3'b111;
        rom_memory[18593] = 3'b110;
        rom_memory[18594] = 3'b111;
        rom_memory[18595] = 3'b111;
        rom_memory[18596] = 3'b111;
        rom_memory[18597] = 3'b110;
        rom_memory[18598] = 3'b110;
        rom_memory[18599] = 3'b110;
        rom_memory[18600] = 3'b110;
        rom_memory[18601] = 3'b110;
        rom_memory[18602] = 3'b110;
        rom_memory[18603] = 3'b110;
        rom_memory[18604] = 3'b110;
        rom_memory[18605] = 3'b110;
        rom_memory[18606] = 3'b110;
        rom_memory[18607] = 3'b110;
        rom_memory[18608] = 3'b110;
        rom_memory[18609] = 3'b110;
        rom_memory[18610] = 3'b110;
        rom_memory[18611] = 3'b110;
        rom_memory[18612] = 3'b110;
        rom_memory[18613] = 3'b111;
        rom_memory[18614] = 3'b110;
        rom_memory[18615] = 3'b110;
        rom_memory[18616] = 3'b110;
        rom_memory[18617] = 3'b110;
        rom_memory[18618] = 3'b110;
        rom_memory[18619] = 3'b110;
        rom_memory[18620] = 3'b110;
        rom_memory[18621] = 3'b111;
        rom_memory[18622] = 3'b111;
        rom_memory[18623] = 3'b111;
        rom_memory[18624] = 3'b111;
        rom_memory[18625] = 3'b111;
        rom_memory[18626] = 3'b111;
        rom_memory[18627] = 3'b111;
        rom_memory[18628] = 3'b111;
        rom_memory[18629] = 3'b111;
        rom_memory[18630] = 3'b111;
        rom_memory[18631] = 3'b111;
        rom_memory[18632] = 3'b111;
        rom_memory[18633] = 3'b111;
        rom_memory[18634] = 3'b111;
        rom_memory[18635] = 3'b111;
        rom_memory[18636] = 3'b111;
        rom_memory[18637] = 3'b111;
        rom_memory[18638] = 3'b111;
        rom_memory[18639] = 3'b111;
        rom_memory[18640] = 3'b111;
        rom_memory[18641] = 3'b111;
        rom_memory[18642] = 3'b111;
        rom_memory[18643] = 3'b111;
        rom_memory[18644] = 3'b111;
        rom_memory[18645] = 3'b111;
        rom_memory[18646] = 3'b111;
        rom_memory[18647] = 3'b111;
        rom_memory[18648] = 3'b111;
        rom_memory[18649] = 3'b111;
        rom_memory[18650] = 3'b111;
        rom_memory[18651] = 3'b111;
        rom_memory[18652] = 3'b111;
        rom_memory[18653] = 3'b111;
        rom_memory[18654] = 3'b111;
        rom_memory[18655] = 3'b111;
        rom_memory[18656] = 3'b111;
        rom_memory[18657] = 3'b111;
        rom_memory[18658] = 3'b111;
        rom_memory[18659] = 3'b111;
        rom_memory[18660] = 3'b111;
        rom_memory[18661] = 3'b111;
        rom_memory[18662] = 3'b111;
        rom_memory[18663] = 3'b111;
        rom_memory[18664] = 3'b111;
        rom_memory[18665] = 3'b111;
        rom_memory[18666] = 3'b110;
        rom_memory[18667] = 3'b110;
        rom_memory[18668] = 3'b110;
        rom_memory[18669] = 3'b111;
        rom_memory[18670] = 3'b111;
        rom_memory[18671] = 3'b110;
        rom_memory[18672] = 3'b110;
        rom_memory[18673] = 3'b110;
        rom_memory[18674] = 3'b110;
        rom_memory[18675] = 3'b110;
        rom_memory[18676] = 3'b110;
        rom_memory[18677] = 3'b110;
        rom_memory[18678] = 3'b110;
        rom_memory[18679] = 3'b110;
        rom_memory[18680] = 3'b110;
        rom_memory[18681] = 3'b110;
        rom_memory[18682] = 3'b110;
        rom_memory[18683] = 3'b110;
        rom_memory[18684] = 3'b110;
        rom_memory[18685] = 3'b110;
        rom_memory[18686] = 3'b110;
        rom_memory[18687] = 3'b110;
        rom_memory[18688] = 3'b110;
        rom_memory[18689] = 3'b110;
        rom_memory[18690] = 3'b110;
        rom_memory[18691] = 3'b110;
        rom_memory[18692] = 3'b110;
        rom_memory[18693] = 3'b110;
        rom_memory[18694] = 3'b110;
        rom_memory[18695] = 3'b110;
        rom_memory[18696] = 3'b110;
        rom_memory[18697] = 3'b110;
        rom_memory[18698] = 3'b110;
        rom_memory[18699] = 3'b110;
        rom_memory[18700] = 3'b110;
        rom_memory[18701] = 3'b110;
        rom_memory[18702] = 3'b110;
        rom_memory[18703] = 3'b110;
        rom_memory[18704] = 3'b110;
        rom_memory[18705] = 3'b110;
        rom_memory[18706] = 3'b110;
        rom_memory[18707] = 3'b110;
        rom_memory[18708] = 3'b110;
        rom_memory[18709] = 3'b110;
        rom_memory[18710] = 3'b110;
        rom_memory[18711] = 3'b110;
        rom_memory[18712] = 3'b110;
        rom_memory[18713] = 3'b110;
        rom_memory[18714] = 3'b110;
        rom_memory[18715] = 3'b110;
        rom_memory[18716] = 3'b110;
        rom_memory[18717] = 3'b110;
        rom_memory[18718] = 3'b110;
        rom_memory[18719] = 3'b110;
        rom_memory[18720] = 3'b110;
        rom_memory[18721] = 3'b110;
        rom_memory[18722] = 3'b110;
        rom_memory[18723] = 3'b110;
        rom_memory[18724] = 3'b110;
        rom_memory[18725] = 3'b110;
        rom_memory[18726] = 3'b110;
        rom_memory[18727] = 3'b110;
        rom_memory[18728] = 3'b110;
        rom_memory[18729] = 3'b110;
        rom_memory[18730] = 3'b110;
        rom_memory[18731] = 3'b110;
        rom_memory[18732] = 3'b110;
        rom_memory[18733] = 3'b110;
        rom_memory[18734] = 3'b110;
        rom_memory[18735] = 3'b110;
        rom_memory[18736] = 3'b110;
        rom_memory[18737] = 3'b110;
        rom_memory[18738] = 3'b110;
        rom_memory[18739] = 3'b110;
        rom_memory[18740] = 3'b110;
        rom_memory[18741] = 3'b110;
        rom_memory[18742] = 3'b110;
        rom_memory[18743] = 3'b110;
        rom_memory[18744] = 3'b110;
        rom_memory[18745] = 3'b110;
        rom_memory[18746] = 3'b110;
        rom_memory[18747] = 3'b110;
        rom_memory[18748] = 3'b110;
        rom_memory[18749] = 3'b110;
        rom_memory[18750] = 3'b111;
        rom_memory[18751] = 3'b111;
        rom_memory[18752] = 3'b111;
        rom_memory[18753] = 3'b111;
        rom_memory[18754] = 3'b111;
        rom_memory[18755] = 3'b111;
        rom_memory[18756] = 3'b111;
        rom_memory[18757] = 3'b111;
        rom_memory[18758] = 3'b111;
        rom_memory[18759] = 3'b111;
        rom_memory[18760] = 3'b111;
        rom_memory[18761] = 3'b111;
        rom_memory[18762] = 3'b111;
        rom_memory[18763] = 3'b111;
        rom_memory[18764] = 3'b111;
        rom_memory[18765] = 3'b110;
        rom_memory[18766] = 3'b100;
        rom_memory[18767] = 3'b100;
        rom_memory[18768] = 3'b100;
        rom_memory[18769] = 3'b100;
        rom_memory[18770] = 3'b110;
        rom_memory[18771] = 3'b110;
        rom_memory[18772] = 3'b110;
        rom_memory[18773] = 3'b110;
        rom_memory[18774] = 3'b100;
        rom_memory[18775] = 3'b110;
        rom_memory[18776] = 3'b100;
        rom_memory[18777] = 3'b110;
        rom_memory[18778] = 3'b110;
        rom_memory[18779] = 3'b100;
        rom_memory[18780] = 3'b100;
        rom_memory[18781] = 3'b100;
        rom_memory[18782] = 3'b100;
        rom_memory[18783] = 3'b100;
        rom_memory[18784] = 3'b110;
        rom_memory[18785] = 3'b110;
        rom_memory[18786] = 3'b110;
        rom_memory[18787] = 3'b110;
        rom_memory[18788] = 3'b110;
        rom_memory[18789] = 3'b110;
        rom_memory[18790] = 3'b110;
        rom_memory[18791] = 3'b110;
        rom_memory[18792] = 3'b110;
        rom_memory[18793] = 3'b110;
        rom_memory[18794] = 3'b110;
        rom_memory[18795] = 3'b110;
        rom_memory[18796] = 3'b110;
        rom_memory[18797] = 3'b110;
        rom_memory[18798] = 3'b110;
        rom_memory[18799] = 3'b110;
        rom_memory[18800] = 3'b110;
        rom_memory[18801] = 3'b110;
        rom_memory[18802] = 3'b110;
        rom_memory[18803] = 3'b110;
        rom_memory[18804] = 3'b110;
        rom_memory[18805] = 3'b110;
        rom_memory[18806] = 3'b110;
        rom_memory[18807] = 3'b110;
        rom_memory[18808] = 3'b110;
        rom_memory[18809] = 3'b110;
        rom_memory[18810] = 3'b110;
        rom_memory[18811] = 3'b110;
        rom_memory[18812] = 3'b110;
        rom_memory[18813] = 3'b110;
        rom_memory[18814] = 3'b100;
        rom_memory[18815] = 3'b000;
        rom_memory[18816] = 3'b000;
        rom_memory[18817] = 3'b000;
        rom_memory[18818] = 3'b000;
        rom_memory[18819] = 3'b000;
        rom_memory[18820] = 3'b100;
        rom_memory[18821] = 3'b100;
        rom_memory[18822] = 3'b100;
        rom_memory[18823] = 3'b110;
        rom_memory[18824] = 3'b110;
        rom_memory[18825] = 3'b110;
        rom_memory[18826] = 3'b000;
        rom_memory[18827] = 3'b000;
        rom_memory[18828] = 3'b110;
        rom_memory[18829] = 3'b100;
        rom_memory[18830] = 3'b000;
        rom_memory[18831] = 3'b110;
        rom_memory[18832] = 3'b111;
        rom_memory[18833] = 3'b111;
        rom_memory[18834] = 3'b110;
        rom_memory[18835] = 3'b110;
        rom_memory[18836] = 3'b110;
        rom_memory[18837] = 3'b111;
        rom_memory[18838] = 3'b110;
        rom_memory[18839] = 3'b110;
        rom_memory[18840] = 3'b110;
        rom_memory[18841] = 3'b110;
        rom_memory[18842] = 3'b110;
        rom_memory[18843] = 3'b110;
        rom_memory[18844] = 3'b110;
        rom_memory[18845] = 3'b110;
        rom_memory[18846] = 3'b110;
        rom_memory[18847] = 3'b110;
        rom_memory[18848] = 3'b110;
        rom_memory[18849] = 3'b110;
        rom_memory[18850] = 3'b110;
        rom_memory[18851] = 3'b110;
        rom_memory[18852] = 3'b110;
        rom_memory[18853] = 3'b110;
        rom_memory[18854] = 3'b110;
        rom_memory[18855] = 3'b110;
        rom_memory[18856] = 3'b110;
        rom_memory[18857] = 3'b110;
        rom_memory[18858] = 3'b110;
        rom_memory[18859] = 3'b110;
        rom_memory[18860] = 3'b111;
        rom_memory[18861] = 3'b111;
        rom_memory[18862] = 3'b111;
        rom_memory[18863] = 3'b111;
        rom_memory[18864] = 3'b111;
        rom_memory[18865] = 3'b111;
        rom_memory[18866] = 3'b111;
        rom_memory[18867] = 3'b111;
        rom_memory[18868] = 3'b111;
        rom_memory[18869] = 3'b111;
        rom_memory[18870] = 3'b111;
        rom_memory[18871] = 3'b111;
        rom_memory[18872] = 3'b111;
        rom_memory[18873] = 3'b111;
        rom_memory[18874] = 3'b111;
        rom_memory[18875] = 3'b111;
        rom_memory[18876] = 3'b111;
        rom_memory[18877] = 3'b111;
        rom_memory[18878] = 3'b111;
        rom_memory[18879] = 3'b111;
        rom_memory[18880] = 3'b111;
        rom_memory[18881] = 3'b111;
        rom_memory[18882] = 3'b111;
        rom_memory[18883] = 3'b111;
        rom_memory[18884] = 3'b111;
        rom_memory[18885] = 3'b111;
        rom_memory[18886] = 3'b111;
        rom_memory[18887] = 3'b111;
        rom_memory[18888] = 3'b111;
        rom_memory[18889] = 3'b111;
        rom_memory[18890] = 3'b111;
        rom_memory[18891] = 3'b111;
        rom_memory[18892] = 3'b111;
        rom_memory[18893] = 3'b111;
        rom_memory[18894] = 3'b111;
        rom_memory[18895] = 3'b111;
        rom_memory[18896] = 3'b111;
        rom_memory[18897] = 3'b111;
        rom_memory[18898] = 3'b111;
        rom_memory[18899] = 3'b111;
        rom_memory[18900] = 3'b111;
        rom_memory[18901] = 3'b111;
        rom_memory[18902] = 3'b111;
        rom_memory[18903] = 3'b111;
        rom_memory[18904] = 3'b111;
        rom_memory[18905] = 3'b111;
        rom_memory[18906] = 3'b110;
        rom_memory[18907] = 3'b110;
        rom_memory[18908] = 3'b110;
        rom_memory[18909] = 3'b111;
        rom_memory[18910] = 3'b110;
        rom_memory[18911] = 3'b110;
        rom_memory[18912] = 3'b110;
        rom_memory[18913] = 3'b110;
        rom_memory[18914] = 3'b110;
        rom_memory[18915] = 3'b110;
        rom_memory[18916] = 3'b110;
        rom_memory[18917] = 3'b110;
        rom_memory[18918] = 3'b110;
        rom_memory[18919] = 3'b110;
        rom_memory[18920] = 3'b110;
        rom_memory[18921] = 3'b110;
        rom_memory[18922] = 3'b110;
        rom_memory[18923] = 3'b110;
        rom_memory[18924] = 3'b110;
        rom_memory[18925] = 3'b110;
        rom_memory[18926] = 3'b110;
        rom_memory[18927] = 3'b110;
        rom_memory[18928] = 3'b110;
        rom_memory[18929] = 3'b110;
        rom_memory[18930] = 3'b110;
        rom_memory[18931] = 3'b110;
        rom_memory[18932] = 3'b110;
        rom_memory[18933] = 3'b110;
        rom_memory[18934] = 3'b110;
        rom_memory[18935] = 3'b110;
        rom_memory[18936] = 3'b110;
        rom_memory[18937] = 3'b110;
        rom_memory[18938] = 3'b110;
        rom_memory[18939] = 3'b110;
        rom_memory[18940] = 3'b110;
        rom_memory[18941] = 3'b110;
        rom_memory[18942] = 3'b110;
        rom_memory[18943] = 3'b110;
        rom_memory[18944] = 3'b110;
        rom_memory[18945] = 3'b110;
        rom_memory[18946] = 3'b110;
        rom_memory[18947] = 3'b110;
        rom_memory[18948] = 3'b110;
        rom_memory[18949] = 3'b110;
        rom_memory[18950] = 3'b110;
        rom_memory[18951] = 3'b110;
        rom_memory[18952] = 3'b110;
        rom_memory[18953] = 3'b110;
        rom_memory[18954] = 3'b110;
        rom_memory[18955] = 3'b110;
        rom_memory[18956] = 3'b110;
        rom_memory[18957] = 3'b110;
        rom_memory[18958] = 3'b110;
        rom_memory[18959] = 3'b110;
        rom_memory[18960] = 3'b110;
        rom_memory[18961] = 3'b110;
        rom_memory[18962] = 3'b110;
        rom_memory[18963] = 3'b110;
        rom_memory[18964] = 3'b110;
        rom_memory[18965] = 3'b110;
        rom_memory[18966] = 3'b110;
        rom_memory[18967] = 3'b110;
        rom_memory[18968] = 3'b110;
        rom_memory[18969] = 3'b110;
        rom_memory[18970] = 3'b110;
        rom_memory[18971] = 3'b110;
        rom_memory[18972] = 3'b110;
        rom_memory[18973] = 3'b110;
        rom_memory[18974] = 3'b110;
        rom_memory[18975] = 3'b110;
        rom_memory[18976] = 3'b110;
        rom_memory[18977] = 3'b110;
        rom_memory[18978] = 3'b110;
        rom_memory[18979] = 3'b110;
        rom_memory[18980] = 3'b110;
        rom_memory[18981] = 3'b110;
        rom_memory[18982] = 3'b110;
        rom_memory[18983] = 3'b110;
        rom_memory[18984] = 3'b110;
        rom_memory[18985] = 3'b110;
        rom_memory[18986] = 3'b110;
        rom_memory[18987] = 3'b110;
        rom_memory[18988] = 3'b110;
        rom_memory[18989] = 3'b111;
        rom_memory[18990] = 3'b111;
        rom_memory[18991] = 3'b111;
        rom_memory[18992] = 3'b111;
        rom_memory[18993] = 3'b111;
        rom_memory[18994] = 3'b111;
        rom_memory[18995] = 3'b111;
        rom_memory[18996] = 3'b111;
        rom_memory[18997] = 3'b111;
        rom_memory[18998] = 3'b111;
        rom_memory[18999] = 3'b111;
        rom_memory[19000] = 3'b111;
        rom_memory[19001] = 3'b111;
        rom_memory[19002] = 3'b111;
        rom_memory[19003] = 3'b111;
        rom_memory[19004] = 3'b111;
        rom_memory[19005] = 3'b111;
        rom_memory[19006] = 3'b100;
        rom_memory[19007] = 3'b100;
        rom_memory[19008] = 3'b100;
        rom_memory[19009] = 3'b100;
        rom_memory[19010] = 3'b110;
        rom_memory[19011] = 3'b110;
        rom_memory[19012] = 3'b110;
        rom_memory[19013] = 3'b110;
        rom_memory[19014] = 3'b110;
        rom_memory[19015] = 3'b110;
        rom_memory[19016] = 3'b110;
        rom_memory[19017] = 3'b110;
        rom_memory[19018] = 3'b110;
        rom_memory[19019] = 3'b100;
        rom_memory[19020] = 3'b100;
        rom_memory[19021] = 3'b100;
        rom_memory[19022] = 3'b100;
        rom_memory[19023] = 3'b100;
        rom_memory[19024] = 3'b110;
        rom_memory[19025] = 3'b110;
        rom_memory[19026] = 3'b110;
        rom_memory[19027] = 3'b110;
        rom_memory[19028] = 3'b100;
        rom_memory[19029] = 3'b100;
        rom_memory[19030] = 3'b110;
        rom_memory[19031] = 3'b110;
        rom_memory[19032] = 3'b110;
        rom_memory[19033] = 3'b100;
        rom_memory[19034] = 3'b110;
        rom_memory[19035] = 3'b110;
        rom_memory[19036] = 3'b110;
        rom_memory[19037] = 3'b110;
        rom_memory[19038] = 3'b110;
        rom_memory[19039] = 3'b110;
        rom_memory[19040] = 3'b110;
        rom_memory[19041] = 3'b110;
        rom_memory[19042] = 3'b110;
        rom_memory[19043] = 3'b110;
        rom_memory[19044] = 3'b110;
        rom_memory[19045] = 3'b110;
        rom_memory[19046] = 3'b110;
        rom_memory[19047] = 3'b110;
        rom_memory[19048] = 3'b110;
        rom_memory[19049] = 3'b110;
        rom_memory[19050] = 3'b110;
        rom_memory[19051] = 3'b110;
        rom_memory[19052] = 3'b110;
        rom_memory[19053] = 3'b100;
        rom_memory[19054] = 3'b110;
        rom_memory[19055] = 3'b110;
        rom_memory[19056] = 3'b000;
        rom_memory[19057] = 3'b000;
        rom_memory[19058] = 3'b000;
        rom_memory[19059] = 3'b000;
        rom_memory[19060] = 3'b000;
        rom_memory[19061] = 3'b100;
        rom_memory[19062] = 3'b000;
        rom_memory[19063] = 3'b100;
        rom_memory[19064] = 3'b110;
        rom_memory[19065] = 3'b110;
        rom_memory[19066] = 3'b100;
        rom_memory[19067] = 3'b000;
        rom_memory[19068] = 3'b000;
        rom_memory[19069] = 3'b110;
        rom_memory[19070] = 3'b100;
        rom_memory[19071] = 3'b000;
        rom_memory[19072] = 3'b100;
        rom_memory[19073] = 3'b110;
        rom_memory[19074] = 3'b110;
        rom_memory[19075] = 3'b110;
        rom_memory[19076] = 3'b110;
        rom_memory[19077] = 3'b110;
        rom_memory[19078] = 3'b111;
        rom_memory[19079] = 3'b110;
        rom_memory[19080] = 3'b110;
        rom_memory[19081] = 3'b110;
        rom_memory[19082] = 3'b110;
        rom_memory[19083] = 3'b110;
        rom_memory[19084] = 3'b110;
        rom_memory[19085] = 3'b110;
        rom_memory[19086] = 3'b110;
        rom_memory[19087] = 3'b110;
        rom_memory[19088] = 3'b110;
        rom_memory[19089] = 3'b110;
        rom_memory[19090] = 3'b110;
        rom_memory[19091] = 3'b110;
        rom_memory[19092] = 3'b110;
        rom_memory[19093] = 3'b110;
        rom_memory[19094] = 3'b110;
        rom_memory[19095] = 3'b110;
        rom_memory[19096] = 3'b111;
        rom_memory[19097] = 3'b110;
        rom_memory[19098] = 3'b110;
        rom_memory[19099] = 3'b111;
        rom_memory[19100] = 3'b110;
        rom_memory[19101] = 3'b110;
        rom_memory[19102] = 3'b111;
        rom_memory[19103] = 3'b111;
        rom_memory[19104] = 3'b111;
        rom_memory[19105] = 3'b111;
        rom_memory[19106] = 3'b111;
        rom_memory[19107] = 3'b111;
        rom_memory[19108] = 3'b111;
        rom_memory[19109] = 3'b111;
        rom_memory[19110] = 3'b111;
        rom_memory[19111] = 3'b111;
        rom_memory[19112] = 3'b111;
        rom_memory[19113] = 3'b111;
        rom_memory[19114] = 3'b111;
        rom_memory[19115] = 3'b111;
        rom_memory[19116] = 3'b111;
        rom_memory[19117] = 3'b111;
        rom_memory[19118] = 3'b111;
        rom_memory[19119] = 3'b111;
        rom_memory[19120] = 3'b111;
        rom_memory[19121] = 3'b111;
        rom_memory[19122] = 3'b111;
        rom_memory[19123] = 3'b111;
        rom_memory[19124] = 3'b111;
        rom_memory[19125] = 3'b111;
        rom_memory[19126] = 3'b111;
        rom_memory[19127] = 3'b111;
        rom_memory[19128] = 3'b111;
        rom_memory[19129] = 3'b111;
        rom_memory[19130] = 3'b111;
        rom_memory[19131] = 3'b111;
        rom_memory[19132] = 3'b111;
        rom_memory[19133] = 3'b111;
        rom_memory[19134] = 3'b111;
        rom_memory[19135] = 3'b111;
        rom_memory[19136] = 3'b111;
        rom_memory[19137] = 3'b111;
        rom_memory[19138] = 3'b111;
        rom_memory[19139] = 3'b111;
        rom_memory[19140] = 3'b111;
        rom_memory[19141] = 3'b111;
        rom_memory[19142] = 3'b111;
        rom_memory[19143] = 3'b111;
        rom_memory[19144] = 3'b111;
        rom_memory[19145] = 3'b111;
        rom_memory[19146] = 3'b110;
        rom_memory[19147] = 3'b110;
        rom_memory[19148] = 3'b110;
        rom_memory[19149] = 3'b110;
        rom_memory[19150] = 3'b111;
        rom_memory[19151] = 3'b110;
        rom_memory[19152] = 3'b110;
        rom_memory[19153] = 3'b110;
        rom_memory[19154] = 3'b110;
        rom_memory[19155] = 3'b110;
        rom_memory[19156] = 3'b110;
        rom_memory[19157] = 3'b110;
        rom_memory[19158] = 3'b110;
        rom_memory[19159] = 3'b110;
        rom_memory[19160] = 3'b110;
        rom_memory[19161] = 3'b110;
        rom_memory[19162] = 3'b110;
        rom_memory[19163] = 3'b110;
        rom_memory[19164] = 3'b110;
        rom_memory[19165] = 3'b110;
        rom_memory[19166] = 3'b110;
        rom_memory[19167] = 3'b110;
        rom_memory[19168] = 3'b110;
        rom_memory[19169] = 3'b110;
        rom_memory[19170] = 3'b110;
        rom_memory[19171] = 3'b110;
        rom_memory[19172] = 3'b110;
        rom_memory[19173] = 3'b110;
        rom_memory[19174] = 3'b110;
        rom_memory[19175] = 3'b110;
        rom_memory[19176] = 3'b110;
        rom_memory[19177] = 3'b110;
        rom_memory[19178] = 3'b110;
        rom_memory[19179] = 3'b110;
        rom_memory[19180] = 3'b110;
        rom_memory[19181] = 3'b110;
        rom_memory[19182] = 3'b110;
        rom_memory[19183] = 3'b110;
        rom_memory[19184] = 3'b110;
        rom_memory[19185] = 3'b110;
        rom_memory[19186] = 3'b110;
        rom_memory[19187] = 3'b110;
        rom_memory[19188] = 3'b110;
        rom_memory[19189] = 3'b110;
        rom_memory[19190] = 3'b110;
        rom_memory[19191] = 3'b110;
        rom_memory[19192] = 3'b110;
        rom_memory[19193] = 3'b110;
        rom_memory[19194] = 3'b110;
        rom_memory[19195] = 3'b110;
        rom_memory[19196] = 3'b110;
        rom_memory[19197] = 3'b110;
        rom_memory[19198] = 3'b110;
        rom_memory[19199] = 3'b110;
        rom_memory[19200] = 3'b110;
        rom_memory[19201] = 3'b110;
        rom_memory[19202] = 3'b110;
        rom_memory[19203] = 3'b110;
        rom_memory[19204] = 3'b110;
        rom_memory[19205] = 3'b110;
        rom_memory[19206] = 3'b110;
        rom_memory[19207] = 3'b110;
        rom_memory[19208] = 3'b110;
        rom_memory[19209] = 3'b110;
        rom_memory[19210] = 3'b110;
        rom_memory[19211] = 3'b110;
        rom_memory[19212] = 3'b110;
        rom_memory[19213] = 3'b110;
        rom_memory[19214] = 3'b110;
        rom_memory[19215] = 3'b110;
        rom_memory[19216] = 3'b110;
        rom_memory[19217] = 3'b110;
        rom_memory[19218] = 3'b110;
        rom_memory[19219] = 3'b110;
        rom_memory[19220] = 3'b110;
        rom_memory[19221] = 3'b110;
        rom_memory[19222] = 3'b110;
        rom_memory[19223] = 3'b110;
        rom_memory[19224] = 3'b110;
        rom_memory[19225] = 3'b110;
        rom_memory[19226] = 3'b110;
        rom_memory[19227] = 3'b110;
        rom_memory[19228] = 3'b110;
        rom_memory[19229] = 3'b111;
        rom_memory[19230] = 3'b111;
        rom_memory[19231] = 3'b111;
        rom_memory[19232] = 3'b111;
        rom_memory[19233] = 3'b111;
        rom_memory[19234] = 3'b111;
        rom_memory[19235] = 3'b111;
        rom_memory[19236] = 3'b111;
        rom_memory[19237] = 3'b111;
        rom_memory[19238] = 3'b111;
        rom_memory[19239] = 3'b111;
        rom_memory[19240] = 3'b111;
        rom_memory[19241] = 3'b111;
        rom_memory[19242] = 3'b111;
        rom_memory[19243] = 3'b111;
        rom_memory[19244] = 3'b111;
        rom_memory[19245] = 3'b111;
        rom_memory[19246] = 3'b110;
        rom_memory[19247] = 3'b100;
        rom_memory[19248] = 3'b100;
        rom_memory[19249] = 3'b100;
        rom_memory[19250] = 3'b110;
        rom_memory[19251] = 3'b110;
        rom_memory[19252] = 3'b110;
        rom_memory[19253] = 3'b110;
        rom_memory[19254] = 3'b110;
        rom_memory[19255] = 3'b110;
        rom_memory[19256] = 3'b100;
        rom_memory[19257] = 3'b100;
        rom_memory[19258] = 3'b110;
        rom_memory[19259] = 3'b110;
        rom_memory[19260] = 3'b110;
        rom_memory[19261] = 3'b100;
        rom_memory[19262] = 3'b100;
        rom_memory[19263] = 3'b100;
        rom_memory[19264] = 3'b110;
        rom_memory[19265] = 3'b110;
        rom_memory[19266] = 3'b110;
        rom_memory[19267] = 3'b110;
        rom_memory[19268] = 3'b110;
        rom_memory[19269] = 3'b110;
        rom_memory[19270] = 3'b110;
        rom_memory[19271] = 3'b110;
        rom_memory[19272] = 3'b110;
        rom_memory[19273] = 3'b110;
        rom_memory[19274] = 3'b110;
        rom_memory[19275] = 3'b110;
        rom_memory[19276] = 3'b110;
        rom_memory[19277] = 3'b110;
        rom_memory[19278] = 3'b110;
        rom_memory[19279] = 3'b110;
        rom_memory[19280] = 3'b110;
        rom_memory[19281] = 3'b110;
        rom_memory[19282] = 3'b110;
        rom_memory[19283] = 3'b110;
        rom_memory[19284] = 3'b110;
        rom_memory[19285] = 3'b110;
        rom_memory[19286] = 3'b110;
        rom_memory[19287] = 3'b110;
        rom_memory[19288] = 3'b110;
        rom_memory[19289] = 3'b110;
        rom_memory[19290] = 3'b110;
        rom_memory[19291] = 3'b110;
        rom_memory[19292] = 3'b111;
        rom_memory[19293] = 3'b111;
        rom_memory[19294] = 3'b000;
        rom_memory[19295] = 3'b000;
        rom_memory[19296] = 3'b110;
        rom_memory[19297] = 3'b000;
        rom_memory[19298] = 3'b000;
        rom_memory[19299] = 3'b000;
        rom_memory[19300] = 3'b000;
        rom_memory[19301] = 3'b000;
        rom_memory[19302] = 3'b000;
        rom_memory[19303] = 3'b000;
        rom_memory[19304] = 3'b100;
        rom_memory[19305] = 3'b110;
        rom_memory[19306] = 3'b110;
        rom_memory[19307] = 3'b000;
        rom_memory[19308] = 3'b000;
        rom_memory[19309] = 3'b000;
        rom_memory[19310] = 3'b110;
        rom_memory[19311] = 3'b110;
        rom_memory[19312] = 3'b110;
        rom_memory[19313] = 3'b110;
        rom_memory[19314] = 3'b110;
        rom_memory[19315] = 3'b110;
        rom_memory[19316] = 3'b110;
        rom_memory[19317] = 3'b110;
        rom_memory[19318] = 3'b111;
        rom_memory[19319] = 3'b111;
        rom_memory[19320] = 3'b110;
        rom_memory[19321] = 3'b110;
        rom_memory[19322] = 3'b110;
        rom_memory[19323] = 3'b110;
        rom_memory[19324] = 3'b110;
        rom_memory[19325] = 3'b110;
        rom_memory[19326] = 3'b110;
        rom_memory[19327] = 3'b110;
        rom_memory[19328] = 3'b110;
        rom_memory[19329] = 3'b110;
        rom_memory[19330] = 3'b110;
        rom_memory[19331] = 3'b110;
        rom_memory[19332] = 3'b110;
        rom_memory[19333] = 3'b110;
        rom_memory[19334] = 3'b110;
        rom_memory[19335] = 3'b110;
        rom_memory[19336] = 3'b110;
        rom_memory[19337] = 3'b110;
        rom_memory[19338] = 3'b110;
        rom_memory[19339] = 3'b111;
        rom_memory[19340] = 3'b110;
        rom_memory[19341] = 3'b111;
        rom_memory[19342] = 3'b111;
        rom_memory[19343] = 3'b111;
        rom_memory[19344] = 3'b111;
        rom_memory[19345] = 3'b111;
        rom_memory[19346] = 3'b111;
        rom_memory[19347] = 3'b111;
        rom_memory[19348] = 3'b111;
        rom_memory[19349] = 3'b111;
        rom_memory[19350] = 3'b111;
        rom_memory[19351] = 3'b111;
        rom_memory[19352] = 3'b111;
        rom_memory[19353] = 3'b111;
        rom_memory[19354] = 3'b111;
        rom_memory[19355] = 3'b111;
        rom_memory[19356] = 3'b111;
        rom_memory[19357] = 3'b111;
        rom_memory[19358] = 3'b111;
        rom_memory[19359] = 3'b111;
        rom_memory[19360] = 3'b111;
        rom_memory[19361] = 3'b111;
        rom_memory[19362] = 3'b111;
        rom_memory[19363] = 3'b111;
        rom_memory[19364] = 3'b111;
        rom_memory[19365] = 3'b111;
        rom_memory[19366] = 3'b111;
        rom_memory[19367] = 3'b111;
        rom_memory[19368] = 3'b111;
        rom_memory[19369] = 3'b111;
        rom_memory[19370] = 3'b111;
        rom_memory[19371] = 3'b111;
        rom_memory[19372] = 3'b111;
        rom_memory[19373] = 3'b111;
        rom_memory[19374] = 3'b111;
        rom_memory[19375] = 3'b111;
        rom_memory[19376] = 3'b111;
        rom_memory[19377] = 3'b111;
        rom_memory[19378] = 3'b111;
        rom_memory[19379] = 3'b111;
        rom_memory[19380] = 3'b111;
        rom_memory[19381] = 3'b111;
        rom_memory[19382] = 3'b111;
        rom_memory[19383] = 3'b111;
        rom_memory[19384] = 3'b111;
        rom_memory[19385] = 3'b111;
        rom_memory[19386] = 3'b110;
        rom_memory[19387] = 3'b110;
        rom_memory[19388] = 3'b110;
        rom_memory[19389] = 3'b111;
        rom_memory[19390] = 3'b111;
        rom_memory[19391] = 3'b111;
        rom_memory[19392] = 3'b110;
        rom_memory[19393] = 3'b110;
        rom_memory[19394] = 3'b110;
        rom_memory[19395] = 3'b110;
        rom_memory[19396] = 3'b110;
        rom_memory[19397] = 3'b110;
        rom_memory[19398] = 3'b110;
        rom_memory[19399] = 3'b110;
        rom_memory[19400] = 3'b110;
        rom_memory[19401] = 3'b110;
        rom_memory[19402] = 3'b110;
        rom_memory[19403] = 3'b110;
        rom_memory[19404] = 3'b110;
        rom_memory[19405] = 3'b110;
        rom_memory[19406] = 3'b110;
        rom_memory[19407] = 3'b110;
        rom_memory[19408] = 3'b110;
        rom_memory[19409] = 3'b110;
        rom_memory[19410] = 3'b110;
        rom_memory[19411] = 3'b110;
        rom_memory[19412] = 3'b110;
        rom_memory[19413] = 3'b110;
        rom_memory[19414] = 3'b110;
        rom_memory[19415] = 3'b110;
        rom_memory[19416] = 3'b110;
        rom_memory[19417] = 3'b110;
        rom_memory[19418] = 3'b110;
        rom_memory[19419] = 3'b110;
        rom_memory[19420] = 3'b110;
        rom_memory[19421] = 3'b110;
        rom_memory[19422] = 3'b110;
        rom_memory[19423] = 3'b110;
        rom_memory[19424] = 3'b110;
        rom_memory[19425] = 3'b110;
        rom_memory[19426] = 3'b110;
        rom_memory[19427] = 3'b110;
        rom_memory[19428] = 3'b110;
        rom_memory[19429] = 3'b110;
        rom_memory[19430] = 3'b110;
        rom_memory[19431] = 3'b110;
        rom_memory[19432] = 3'b110;
        rom_memory[19433] = 3'b110;
        rom_memory[19434] = 3'b110;
        rom_memory[19435] = 3'b110;
        rom_memory[19436] = 3'b110;
        rom_memory[19437] = 3'b110;
        rom_memory[19438] = 3'b110;
        rom_memory[19439] = 3'b110;
        rom_memory[19440] = 3'b110;
        rom_memory[19441] = 3'b110;
        rom_memory[19442] = 3'b110;
        rom_memory[19443] = 3'b110;
        rom_memory[19444] = 3'b110;
        rom_memory[19445] = 3'b110;
        rom_memory[19446] = 3'b110;
        rom_memory[19447] = 3'b110;
        rom_memory[19448] = 3'b110;
        rom_memory[19449] = 3'b110;
        rom_memory[19450] = 3'b110;
        rom_memory[19451] = 3'b110;
        rom_memory[19452] = 3'b110;
        rom_memory[19453] = 3'b110;
        rom_memory[19454] = 3'b110;
        rom_memory[19455] = 3'b110;
        rom_memory[19456] = 3'b110;
        rom_memory[19457] = 3'b110;
        rom_memory[19458] = 3'b110;
        rom_memory[19459] = 3'b110;
        rom_memory[19460] = 3'b110;
        rom_memory[19461] = 3'b110;
        rom_memory[19462] = 3'b110;
        rom_memory[19463] = 3'b110;
        rom_memory[19464] = 3'b110;
        rom_memory[19465] = 3'b110;
        rom_memory[19466] = 3'b110;
        rom_memory[19467] = 3'b110;
        rom_memory[19468] = 3'b110;
        rom_memory[19469] = 3'b111;
        rom_memory[19470] = 3'b111;
        rom_memory[19471] = 3'b111;
        rom_memory[19472] = 3'b111;
        rom_memory[19473] = 3'b111;
        rom_memory[19474] = 3'b111;
        rom_memory[19475] = 3'b111;
        rom_memory[19476] = 3'b111;
        rom_memory[19477] = 3'b111;
        rom_memory[19478] = 3'b111;
        rom_memory[19479] = 3'b111;
        rom_memory[19480] = 3'b111;
        rom_memory[19481] = 3'b111;
        rom_memory[19482] = 3'b111;
        rom_memory[19483] = 3'b111;
        rom_memory[19484] = 3'b111;
        rom_memory[19485] = 3'b111;
        rom_memory[19486] = 3'b110;
        rom_memory[19487] = 3'b100;
        rom_memory[19488] = 3'b100;
        rom_memory[19489] = 3'b100;
        rom_memory[19490] = 3'b110;
        rom_memory[19491] = 3'b110;
        rom_memory[19492] = 3'b100;
        rom_memory[19493] = 3'b110;
        rom_memory[19494] = 3'b110;
        rom_memory[19495] = 3'b110;
        rom_memory[19496] = 3'b110;
        rom_memory[19497] = 3'b100;
        rom_memory[19498] = 3'b110;
        rom_memory[19499] = 3'b110;
        rom_memory[19500] = 3'b110;
        rom_memory[19501] = 3'b110;
        rom_memory[19502] = 3'b100;
        rom_memory[19503] = 3'b100;
        rom_memory[19504] = 3'b100;
        rom_memory[19505] = 3'b110;
        rom_memory[19506] = 3'b110;
        rom_memory[19507] = 3'b110;
        rom_memory[19508] = 3'b110;
        rom_memory[19509] = 3'b110;
        rom_memory[19510] = 3'b110;
        rom_memory[19511] = 3'b110;
        rom_memory[19512] = 3'b110;
        rom_memory[19513] = 3'b110;
        rom_memory[19514] = 3'b110;
        rom_memory[19515] = 3'b110;
        rom_memory[19516] = 3'b110;
        rom_memory[19517] = 3'b110;
        rom_memory[19518] = 3'b110;
        rom_memory[19519] = 3'b110;
        rom_memory[19520] = 3'b110;
        rom_memory[19521] = 3'b110;
        rom_memory[19522] = 3'b110;
        rom_memory[19523] = 3'b110;
        rom_memory[19524] = 3'b110;
        rom_memory[19525] = 3'b110;
        rom_memory[19526] = 3'b110;
        rom_memory[19527] = 3'b110;
        rom_memory[19528] = 3'b110;
        rom_memory[19529] = 3'b110;
        rom_memory[19530] = 3'b110;
        rom_memory[19531] = 3'b110;
        rom_memory[19532] = 3'b110;
        rom_memory[19533] = 3'b111;
        rom_memory[19534] = 3'b111;
        rom_memory[19535] = 3'b000;
        rom_memory[19536] = 3'b000;
        rom_memory[19537] = 3'b000;
        rom_memory[19538] = 3'b000;
        rom_memory[19539] = 3'b000;
        rom_memory[19540] = 3'b000;
        rom_memory[19541] = 3'b000;
        rom_memory[19542] = 3'b000;
        rom_memory[19543] = 3'b000;
        rom_memory[19544] = 3'b000;
        rom_memory[19545] = 3'b110;
        rom_memory[19546] = 3'b110;
        rom_memory[19547] = 3'b110;
        rom_memory[19548] = 3'b000;
        rom_memory[19549] = 3'b000;
        rom_memory[19550] = 3'b100;
        rom_memory[19551] = 3'b110;
        rom_memory[19552] = 3'b110;
        rom_memory[19553] = 3'b110;
        rom_memory[19554] = 3'b110;
        rom_memory[19555] = 3'b110;
        rom_memory[19556] = 3'b110;
        rom_memory[19557] = 3'b110;
        rom_memory[19558] = 3'b111;
        rom_memory[19559] = 3'b111;
        rom_memory[19560] = 3'b111;
        rom_memory[19561] = 3'b110;
        rom_memory[19562] = 3'b110;
        rom_memory[19563] = 3'b110;
        rom_memory[19564] = 3'b110;
        rom_memory[19565] = 3'b110;
        rom_memory[19566] = 3'b110;
        rom_memory[19567] = 3'b110;
        rom_memory[19568] = 3'b110;
        rom_memory[19569] = 3'b110;
        rom_memory[19570] = 3'b110;
        rom_memory[19571] = 3'b110;
        rom_memory[19572] = 3'b110;
        rom_memory[19573] = 3'b110;
        rom_memory[19574] = 3'b110;
        rom_memory[19575] = 3'b110;
        rom_memory[19576] = 3'b110;
        rom_memory[19577] = 3'b110;
        rom_memory[19578] = 3'b110;
        rom_memory[19579] = 3'b110;
        rom_memory[19580] = 3'b110;
        rom_memory[19581] = 3'b111;
        rom_memory[19582] = 3'b111;
        rom_memory[19583] = 3'b111;
        rom_memory[19584] = 3'b111;
        rom_memory[19585] = 3'b111;
        rom_memory[19586] = 3'b111;
        rom_memory[19587] = 3'b111;
        rom_memory[19588] = 3'b111;
        rom_memory[19589] = 3'b111;
        rom_memory[19590] = 3'b111;
        rom_memory[19591] = 3'b111;
        rom_memory[19592] = 3'b111;
        rom_memory[19593] = 3'b111;
        rom_memory[19594] = 3'b111;
        rom_memory[19595] = 3'b111;
        rom_memory[19596] = 3'b111;
        rom_memory[19597] = 3'b111;
        rom_memory[19598] = 3'b111;
        rom_memory[19599] = 3'b111;
        rom_memory[19600] = 3'b111;
        rom_memory[19601] = 3'b111;
        rom_memory[19602] = 3'b111;
        rom_memory[19603] = 3'b111;
        rom_memory[19604] = 3'b111;
        rom_memory[19605] = 3'b111;
        rom_memory[19606] = 3'b111;
        rom_memory[19607] = 3'b111;
        rom_memory[19608] = 3'b111;
        rom_memory[19609] = 3'b111;
        rom_memory[19610] = 3'b111;
        rom_memory[19611] = 3'b111;
        rom_memory[19612] = 3'b111;
        rom_memory[19613] = 3'b111;
        rom_memory[19614] = 3'b111;
        rom_memory[19615] = 3'b111;
        rom_memory[19616] = 3'b111;
        rom_memory[19617] = 3'b111;
        rom_memory[19618] = 3'b111;
        rom_memory[19619] = 3'b111;
        rom_memory[19620] = 3'b111;
        rom_memory[19621] = 3'b111;
        rom_memory[19622] = 3'b111;
        rom_memory[19623] = 3'b111;
        rom_memory[19624] = 3'b111;
        rom_memory[19625] = 3'b110;
        rom_memory[19626] = 3'b111;
        rom_memory[19627] = 3'b111;
        rom_memory[19628] = 3'b111;
        rom_memory[19629] = 3'b110;
        rom_memory[19630] = 3'b110;
        rom_memory[19631] = 3'b111;
        rom_memory[19632] = 3'b110;
        rom_memory[19633] = 3'b110;
        rom_memory[19634] = 3'b110;
        rom_memory[19635] = 3'b110;
        rom_memory[19636] = 3'b110;
        rom_memory[19637] = 3'b110;
        rom_memory[19638] = 3'b110;
        rom_memory[19639] = 3'b110;
        rom_memory[19640] = 3'b110;
        rom_memory[19641] = 3'b110;
        rom_memory[19642] = 3'b110;
        rom_memory[19643] = 3'b110;
        rom_memory[19644] = 3'b110;
        rom_memory[19645] = 3'b110;
        rom_memory[19646] = 3'b110;
        rom_memory[19647] = 3'b110;
        rom_memory[19648] = 3'b110;
        rom_memory[19649] = 3'b110;
        rom_memory[19650] = 3'b110;
        rom_memory[19651] = 3'b110;
        rom_memory[19652] = 3'b110;
        rom_memory[19653] = 3'b110;
        rom_memory[19654] = 3'b110;
        rom_memory[19655] = 3'b110;
        rom_memory[19656] = 3'b110;
        rom_memory[19657] = 3'b110;
        rom_memory[19658] = 3'b110;
        rom_memory[19659] = 3'b110;
        rom_memory[19660] = 3'b110;
        rom_memory[19661] = 3'b110;
        rom_memory[19662] = 3'b110;
        rom_memory[19663] = 3'b110;
        rom_memory[19664] = 3'b110;
        rom_memory[19665] = 3'b110;
        rom_memory[19666] = 3'b110;
        rom_memory[19667] = 3'b110;
        rom_memory[19668] = 3'b110;
        rom_memory[19669] = 3'b110;
        rom_memory[19670] = 3'b110;
        rom_memory[19671] = 3'b110;
        rom_memory[19672] = 3'b110;
        rom_memory[19673] = 3'b110;
        rom_memory[19674] = 3'b110;
        rom_memory[19675] = 3'b110;
        rom_memory[19676] = 3'b110;
        rom_memory[19677] = 3'b110;
        rom_memory[19678] = 3'b110;
        rom_memory[19679] = 3'b110;
        rom_memory[19680] = 3'b110;
        rom_memory[19681] = 3'b110;
        rom_memory[19682] = 3'b110;
        rom_memory[19683] = 3'b110;
        rom_memory[19684] = 3'b110;
        rom_memory[19685] = 3'b110;
        rom_memory[19686] = 3'b110;
        rom_memory[19687] = 3'b110;
        rom_memory[19688] = 3'b110;
        rom_memory[19689] = 3'b110;
        rom_memory[19690] = 3'b110;
        rom_memory[19691] = 3'b110;
        rom_memory[19692] = 3'b110;
        rom_memory[19693] = 3'b110;
        rom_memory[19694] = 3'b110;
        rom_memory[19695] = 3'b110;
        rom_memory[19696] = 3'b110;
        rom_memory[19697] = 3'b110;
        rom_memory[19698] = 3'b110;
        rom_memory[19699] = 3'b110;
        rom_memory[19700] = 3'b110;
        rom_memory[19701] = 3'b110;
        rom_memory[19702] = 3'b110;
        rom_memory[19703] = 3'b110;
        rom_memory[19704] = 3'b110;
        rom_memory[19705] = 3'b110;
        rom_memory[19706] = 3'b110;
        rom_memory[19707] = 3'b110;
        rom_memory[19708] = 3'b110;
        rom_memory[19709] = 3'b110;
        rom_memory[19710] = 3'b111;
        rom_memory[19711] = 3'b111;
        rom_memory[19712] = 3'b111;
        rom_memory[19713] = 3'b111;
        rom_memory[19714] = 3'b111;
        rom_memory[19715] = 3'b111;
        rom_memory[19716] = 3'b111;
        rom_memory[19717] = 3'b111;
        rom_memory[19718] = 3'b111;
        rom_memory[19719] = 3'b111;
        rom_memory[19720] = 3'b111;
        rom_memory[19721] = 3'b111;
        rom_memory[19722] = 3'b111;
        rom_memory[19723] = 3'b111;
        rom_memory[19724] = 3'b111;
        rom_memory[19725] = 3'b111;
        rom_memory[19726] = 3'b110;
        rom_memory[19727] = 3'b100;
        rom_memory[19728] = 3'b100;
        rom_memory[19729] = 3'b100;
        rom_memory[19730] = 3'b110;
        rom_memory[19731] = 3'b110;
        rom_memory[19732] = 3'b100;
        rom_memory[19733] = 3'b110;
        rom_memory[19734] = 3'b110;
        rom_memory[19735] = 3'b110;
        rom_memory[19736] = 3'b110;
        rom_memory[19737] = 3'b100;
        rom_memory[19738] = 3'b110;
        rom_memory[19739] = 3'b110;
        rom_memory[19740] = 3'b110;
        rom_memory[19741] = 3'b110;
        rom_memory[19742] = 3'b110;
        rom_memory[19743] = 3'b100;
        rom_memory[19744] = 3'b100;
        rom_memory[19745] = 3'b100;
        rom_memory[19746] = 3'b110;
        rom_memory[19747] = 3'b110;
        rom_memory[19748] = 3'b110;
        rom_memory[19749] = 3'b110;
        rom_memory[19750] = 3'b110;
        rom_memory[19751] = 3'b110;
        rom_memory[19752] = 3'b110;
        rom_memory[19753] = 3'b110;
        rom_memory[19754] = 3'b110;
        rom_memory[19755] = 3'b110;
        rom_memory[19756] = 3'b110;
        rom_memory[19757] = 3'b110;
        rom_memory[19758] = 3'b110;
        rom_memory[19759] = 3'b110;
        rom_memory[19760] = 3'b110;
        rom_memory[19761] = 3'b110;
        rom_memory[19762] = 3'b110;
        rom_memory[19763] = 3'b100;
        rom_memory[19764] = 3'b110;
        rom_memory[19765] = 3'b110;
        rom_memory[19766] = 3'b110;
        rom_memory[19767] = 3'b110;
        rom_memory[19768] = 3'b110;
        rom_memory[19769] = 3'b110;
        rom_memory[19770] = 3'b110;
        rom_memory[19771] = 3'b110;
        rom_memory[19772] = 3'b110;
        rom_memory[19773] = 3'b110;
        rom_memory[19774] = 3'b111;
        rom_memory[19775] = 3'b111;
        rom_memory[19776] = 3'b000;
        rom_memory[19777] = 3'b000;
        rom_memory[19778] = 3'b000;
        rom_memory[19779] = 3'b000;
        rom_memory[19780] = 3'b000;
        rom_memory[19781] = 3'b000;
        rom_memory[19782] = 3'b000;
        rom_memory[19783] = 3'b000;
        rom_memory[19784] = 3'b000;
        rom_memory[19785] = 3'b100;
        rom_memory[19786] = 3'b110;
        rom_memory[19787] = 3'b110;
        rom_memory[19788] = 3'b110;
        rom_memory[19789] = 3'b100;
        rom_memory[19790] = 3'b110;
        rom_memory[19791] = 3'b110;
        rom_memory[19792] = 3'b110;
        rom_memory[19793] = 3'b110;
        rom_memory[19794] = 3'b110;
        rom_memory[19795] = 3'b110;
        rom_memory[19796] = 3'b110;
        rom_memory[19797] = 3'b110;
        rom_memory[19798] = 3'b110;
        rom_memory[19799] = 3'b111;
        rom_memory[19800] = 3'b111;
        rom_memory[19801] = 3'b111;
        rom_memory[19802] = 3'b110;
        rom_memory[19803] = 3'b110;
        rom_memory[19804] = 3'b110;
        rom_memory[19805] = 3'b110;
        rom_memory[19806] = 3'b110;
        rom_memory[19807] = 3'b110;
        rom_memory[19808] = 3'b110;
        rom_memory[19809] = 3'b110;
        rom_memory[19810] = 3'b110;
        rom_memory[19811] = 3'b110;
        rom_memory[19812] = 3'b110;
        rom_memory[19813] = 3'b110;
        rom_memory[19814] = 3'b110;
        rom_memory[19815] = 3'b110;
        rom_memory[19816] = 3'b110;
        rom_memory[19817] = 3'b110;
        rom_memory[19818] = 3'b110;
        rom_memory[19819] = 3'b110;
        rom_memory[19820] = 3'b111;
        rom_memory[19821] = 3'b111;
        rom_memory[19822] = 3'b111;
        rom_memory[19823] = 3'b111;
        rom_memory[19824] = 3'b111;
        rom_memory[19825] = 3'b111;
        rom_memory[19826] = 3'b111;
        rom_memory[19827] = 3'b111;
        rom_memory[19828] = 3'b111;
        rom_memory[19829] = 3'b111;
        rom_memory[19830] = 3'b111;
        rom_memory[19831] = 3'b111;
        rom_memory[19832] = 3'b111;
        rom_memory[19833] = 3'b111;
        rom_memory[19834] = 3'b111;
        rom_memory[19835] = 3'b111;
        rom_memory[19836] = 3'b111;
        rom_memory[19837] = 3'b111;
        rom_memory[19838] = 3'b111;
        rom_memory[19839] = 3'b111;
        rom_memory[19840] = 3'b111;
        rom_memory[19841] = 3'b111;
        rom_memory[19842] = 3'b111;
        rom_memory[19843] = 3'b111;
        rom_memory[19844] = 3'b111;
        rom_memory[19845] = 3'b111;
        rom_memory[19846] = 3'b111;
        rom_memory[19847] = 3'b111;
        rom_memory[19848] = 3'b111;
        rom_memory[19849] = 3'b111;
        rom_memory[19850] = 3'b111;
        rom_memory[19851] = 3'b111;
        rom_memory[19852] = 3'b111;
        rom_memory[19853] = 3'b111;
        rom_memory[19854] = 3'b111;
        rom_memory[19855] = 3'b111;
        rom_memory[19856] = 3'b111;
        rom_memory[19857] = 3'b111;
        rom_memory[19858] = 3'b111;
        rom_memory[19859] = 3'b111;
        rom_memory[19860] = 3'b111;
        rom_memory[19861] = 3'b111;
        rom_memory[19862] = 3'b111;
        rom_memory[19863] = 3'b111;
        rom_memory[19864] = 3'b111;
        rom_memory[19865] = 3'b111;
        rom_memory[19866] = 3'b110;
        rom_memory[19867] = 3'b111;
        rom_memory[19868] = 3'b111;
        rom_memory[19869] = 3'b111;
        rom_memory[19870] = 3'b110;
        rom_memory[19871] = 3'b110;
        rom_memory[19872] = 3'b110;
        rom_memory[19873] = 3'b110;
        rom_memory[19874] = 3'b110;
        rom_memory[19875] = 3'b110;
        rom_memory[19876] = 3'b110;
        rom_memory[19877] = 3'b110;
        rom_memory[19878] = 3'b110;
        rom_memory[19879] = 3'b110;
        rom_memory[19880] = 3'b110;
        rom_memory[19881] = 3'b110;
        rom_memory[19882] = 3'b110;
        rom_memory[19883] = 3'b110;
        rom_memory[19884] = 3'b110;
        rom_memory[19885] = 3'b110;
        rom_memory[19886] = 3'b110;
        rom_memory[19887] = 3'b110;
        rom_memory[19888] = 3'b110;
        rom_memory[19889] = 3'b110;
        rom_memory[19890] = 3'b110;
        rom_memory[19891] = 3'b110;
        rom_memory[19892] = 3'b110;
        rom_memory[19893] = 3'b110;
        rom_memory[19894] = 3'b110;
        rom_memory[19895] = 3'b110;
        rom_memory[19896] = 3'b110;
        rom_memory[19897] = 3'b110;
        rom_memory[19898] = 3'b110;
        rom_memory[19899] = 3'b110;
        rom_memory[19900] = 3'b110;
        rom_memory[19901] = 3'b110;
        rom_memory[19902] = 3'b110;
        rom_memory[19903] = 3'b110;
        rom_memory[19904] = 3'b110;
        rom_memory[19905] = 3'b110;
        rom_memory[19906] = 3'b110;
        rom_memory[19907] = 3'b110;
        rom_memory[19908] = 3'b110;
        rom_memory[19909] = 3'b110;
        rom_memory[19910] = 3'b110;
        rom_memory[19911] = 3'b110;
        rom_memory[19912] = 3'b110;
        rom_memory[19913] = 3'b110;
        rom_memory[19914] = 3'b110;
        rom_memory[19915] = 3'b110;
        rom_memory[19916] = 3'b110;
        rom_memory[19917] = 3'b110;
        rom_memory[19918] = 3'b110;
        rom_memory[19919] = 3'b110;
        rom_memory[19920] = 3'b110;
        rom_memory[19921] = 3'b110;
        rom_memory[19922] = 3'b110;
        rom_memory[19923] = 3'b110;
        rom_memory[19924] = 3'b110;
        rom_memory[19925] = 3'b110;
        rom_memory[19926] = 3'b110;
        rom_memory[19927] = 3'b110;
        rom_memory[19928] = 3'b110;
        rom_memory[19929] = 3'b110;
        rom_memory[19930] = 3'b110;
        rom_memory[19931] = 3'b110;
        rom_memory[19932] = 3'b110;
        rom_memory[19933] = 3'b110;
        rom_memory[19934] = 3'b110;
        rom_memory[19935] = 3'b110;
        rom_memory[19936] = 3'b110;
        rom_memory[19937] = 3'b110;
        rom_memory[19938] = 3'b110;
        rom_memory[19939] = 3'b110;
        rom_memory[19940] = 3'b110;
        rom_memory[19941] = 3'b110;
        rom_memory[19942] = 3'b110;
        rom_memory[19943] = 3'b110;
        rom_memory[19944] = 3'b110;
        rom_memory[19945] = 3'b110;
        rom_memory[19946] = 3'b110;
        rom_memory[19947] = 3'b110;
        rom_memory[19948] = 3'b110;
        rom_memory[19949] = 3'b110;
        rom_memory[19950] = 3'b111;
        rom_memory[19951] = 3'b111;
        rom_memory[19952] = 3'b111;
        rom_memory[19953] = 3'b111;
        rom_memory[19954] = 3'b111;
        rom_memory[19955] = 3'b111;
        rom_memory[19956] = 3'b111;
        rom_memory[19957] = 3'b111;
        rom_memory[19958] = 3'b111;
        rom_memory[19959] = 3'b111;
        rom_memory[19960] = 3'b111;
        rom_memory[19961] = 3'b111;
        rom_memory[19962] = 3'b111;
        rom_memory[19963] = 3'b111;
        rom_memory[19964] = 3'b111;
        rom_memory[19965] = 3'b111;
        rom_memory[19966] = 3'b110;
        rom_memory[19967] = 3'b100;
        rom_memory[19968] = 3'b100;
        rom_memory[19969] = 3'b100;
        rom_memory[19970] = 3'b110;
        rom_memory[19971] = 3'b110;
        rom_memory[19972] = 3'b110;
        rom_memory[19973] = 3'b110;
        rom_memory[19974] = 3'b110;
        rom_memory[19975] = 3'b110;
        rom_memory[19976] = 3'b110;
        rom_memory[19977] = 3'b110;
        rom_memory[19978] = 3'b110;
        rom_memory[19979] = 3'b110;
        rom_memory[19980] = 3'b110;
        rom_memory[19981] = 3'b110;
        rom_memory[19982] = 3'b110;
        rom_memory[19983] = 3'b100;
        rom_memory[19984] = 3'b100;
        rom_memory[19985] = 3'b100;
        rom_memory[19986] = 3'b100;
        rom_memory[19987] = 3'b110;
        rom_memory[19988] = 3'b110;
        rom_memory[19989] = 3'b110;
        rom_memory[19990] = 3'b110;
        rom_memory[19991] = 3'b110;
        rom_memory[19992] = 3'b110;
        rom_memory[19993] = 3'b110;
        rom_memory[19994] = 3'b110;
        rom_memory[19995] = 3'b110;
        rom_memory[19996] = 3'b110;
        rom_memory[19997] = 3'b110;
        rom_memory[19998] = 3'b110;
        rom_memory[19999] = 3'b110;
        rom_memory[20000] = 3'b110;
        rom_memory[20001] = 3'b110;
        rom_memory[20002] = 3'b110;
        rom_memory[20003] = 3'b110;
        rom_memory[20004] = 3'b110;
        rom_memory[20005] = 3'b110;
        rom_memory[20006] = 3'b110;
        rom_memory[20007] = 3'b110;
        rom_memory[20008] = 3'b110;
        rom_memory[20009] = 3'b110;
        rom_memory[20010] = 3'b110;
        rom_memory[20011] = 3'b110;
        rom_memory[20012] = 3'b110;
        rom_memory[20013] = 3'b110;
        rom_memory[20014] = 3'b110;
        rom_memory[20015] = 3'b111;
        rom_memory[20016] = 3'b000;
        rom_memory[20017] = 3'b000;
        rom_memory[20018] = 3'b000;
        rom_memory[20019] = 3'b000;
        rom_memory[20020] = 3'b000;
        rom_memory[20021] = 3'b000;
        rom_memory[20022] = 3'b000;
        rom_memory[20023] = 3'b000;
        rom_memory[20024] = 3'b000;
        rom_memory[20025] = 3'b000;
        rom_memory[20026] = 3'b000;
        rom_memory[20027] = 3'b000;
        rom_memory[20028] = 3'b000;
        rom_memory[20029] = 3'b000;
        rom_memory[20030] = 3'b000;
        rom_memory[20031] = 3'b110;
        rom_memory[20032] = 3'b110;
        rom_memory[20033] = 3'b110;
        rom_memory[20034] = 3'b110;
        rom_memory[20035] = 3'b110;
        rom_memory[20036] = 3'b110;
        rom_memory[20037] = 3'b110;
        rom_memory[20038] = 3'b110;
        rom_memory[20039] = 3'b110;
        rom_memory[20040] = 3'b111;
        rom_memory[20041] = 3'b111;
        rom_memory[20042] = 3'b111;
        rom_memory[20043] = 3'b110;
        rom_memory[20044] = 3'b110;
        rom_memory[20045] = 3'b110;
        rom_memory[20046] = 3'b110;
        rom_memory[20047] = 3'b110;
        rom_memory[20048] = 3'b110;
        rom_memory[20049] = 3'b110;
        rom_memory[20050] = 3'b110;
        rom_memory[20051] = 3'b110;
        rom_memory[20052] = 3'b110;
        rom_memory[20053] = 3'b110;
        rom_memory[20054] = 3'b110;
        rom_memory[20055] = 3'b110;
        rom_memory[20056] = 3'b110;
        rom_memory[20057] = 3'b110;
        rom_memory[20058] = 3'b110;
        rom_memory[20059] = 3'b110;
        rom_memory[20060] = 3'b111;
        rom_memory[20061] = 3'b110;
        rom_memory[20062] = 3'b111;
        rom_memory[20063] = 3'b111;
        rom_memory[20064] = 3'b111;
        rom_memory[20065] = 3'b111;
        rom_memory[20066] = 3'b111;
        rom_memory[20067] = 3'b111;
        rom_memory[20068] = 3'b111;
        rom_memory[20069] = 3'b111;
        rom_memory[20070] = 3'b111;
        rom_memory[20071] = 3'b111;
        rom_memory[20072] = 3'b111;
        rom_memory[20073] = 3'b111;
        rom_memory[20074] = 3'b111;
        rom_memory[20075] = 3'b111;
        rom_memory[20076] = 3'b111;
        rom_memory[20077] = 3'b111;
        rom_memory[20078] = 3'b111;
        rom_memory[20079] = 3'b111;
        rom_memory[20080] = 3'b111;
        rom_memory[20081] = 3'b111;
        rom_memory[20082] = 3'b111;
        rom_memory[20083] = 3'b111;
        rom_memory[20084] = 3'b111;
        rom_memory[20085] = 3'b111;
        rom_memory[20086] = 3'b111;
        rom_memory[20087] = 3'b111;
        rom_memory[20088] = 3'b111;
        rom_memory[20089] = 3'b111;
        rom_memory[20090] = 3'b111;
        rom_memory[20091] = 3'b111;
        rom_memory[20092] = 3'b111;
        rom_memory[20093] = 3'b111;
        rom_memory[20094] = 3'b111;
        rom_memory[20095] = 3'b111;
        rom_memory[20096] = 3'b111;
        rom_memory[20097] = 3'b111;
        rom_memory[20098] = 3'b111;
        rom_memory[20099] = 3'b111;
        rom_memory[20100] = 3'b111;
        rom_memory[20101] = 3'b111;
        rom_memory[20102] = 3'b111;
        rom_memory[20103] = 3'b111;
        rom_memory[20104] = 3'b111;
        rom_memory[20105] = 3'b111;
        rom_memory[20106] = 3'b111;
        rom_memory[20107] = 3'b111;
        rom_memory[20108] = 3'b111;
        rom_memory[20109] = 3'b110;
        rom_memory[20110] = 3'b110;
        rom_memory[20111] = 3'b110;
        rom_memory[20112] = 3'b110;
        rom_memory[20113] = 3'b110;
        rom_memory[20114] = 3'b110;
        rom_memory[20115] = 3'b110;
        rom_memory[20116] = 3'b110;
        rom_memory[20117] = 3'b110;
        rom_memory[20118] = 3'b110;
        rom_memory[20119] = 3'b110;
        rom_memory[20120] = 3'b110;
        rom_memory[20121] = 3'b110;
        rom_memory[20122] = 3'b110;
        rom_memory[20123] = 3'b110;
        rom_memory[20124] = 3'b110;
        rom_memory[20125] = 3'b110;
        rom_memory[20126] = 3'b110;
        rom_memory[20127] = 3'b110;
        rom_memory[20128] = 3'b110;
        rom_memory[20129] = 3'b110;
        rom_memory[20130] = 3'b110;
        rom_memory[20131] = 3'b110;
        rom_memory[20132] = 3'b110;
        rom_memory[20133] = 3'b110;
        rom_memory[20134] = 3'b110;
        rom_memory[20135] = 3'b110;
        rom_memory[20136] = 3'b110;
        rom_memory[20137] = 3'b110;
        rom_memory[20138] = 3'b110;
        rom_memory[20139] = 3'b110;
        rom_memory[20140] = 3'b110;
        rom_memory[20141] = 3'b110;
        rom_memory[20142] = 3'b110;
        rom_memory[20143] = 3'b110;
        rom_memory[20144] = 3'b110;
        rom_memory[20145] = 3'b110;
        rom_memory[20146] = 3'b110;
        rom_memory[20147] = 3'b110;
        rom_memory[20148] = 3'b110;
        rom_memory[20149] = 3'b110;
        rom_memory[20150] = 3'b110;
        rom_memory[20151] = 3'b110;
        rom_memory[20152] = 3'b110;
        rom_memory[20153] = 3'b110;
        rom_memory[20154] = 3'b110;
        rom_memory[20155] = 3'b110;
        rom_memory[20156] = 3'b110;
        rom_memory[20157] = 3'b110;
        rom_memory[20158] = 3'b110;
        rom_memory[20159] = 3'b110;
        rom_memory[20160] = 3'b110;
        rom_memory[20161] = 3'b110;
        rom_memory[20162] = 3'b110;
        rom_memory[20163] = 3'b110;
        rom_memory[20164] = 3'b110;
        rom_memory[20165] = 3'b110;
        rom_memory[20166] = 3'b110;
        rom_memory[20167] = 3'b110;
        rom_memory[20168] = 3'b110;
        rom_memory[20169] = 3'b110;
        rom_memory[20170] = 3'b110;
        rom_memory[20171] = 3'b110;
        rom_memory[20172] = 3'b110;
        rom_memory[20173] = 3'b110;
        rom_memory[20174] = 3'b110;
        rom_memory[20175] = 3'b110;
        rom_memory[20176] = 3'b110;
        rom_memory[20177] = 3'b110;
        rom_memory[20178] = 3'b110;
        rom_memory[20179] = 3'b110;
        rom_memory[20180] = 3'b110;
        rom_memory[20181] = 3'b110;
        rom_memory[20182] = 3'b110;
        rom_memory[20183] = 3'b110;
        rom_memory[20184] = 3'b110;
        rom_memory[20185] = 3'b110;
        rom_memory[20186] = 3'b110;
        rom_memory[20187] = 3'b110;
        rom_memory[20188] = 3'b110;
        rom_memory[20189] = 3'b110;
        rom_memory[20190] = 3'b111;
        rom_memory[20191] = 3'b111;
        rom_memory[20192] = 3'b111;
        rom_memory[20193] = 3'b111;
        rom_memory[20194] = 3'b111;
        rom_memory[20195] = 3'b111;
        rom_memory[20196] = 3'b111;
        rom_memory[20197] = 3'b111;
        rom_memory[20198] = 3'b111;
        rom_memory[20199] = 3'b111;
        rom_memory[20200] = 3'b111;
        rom_memory[20201] = 3'b111;
        rom_memory[20202] = 3'b111;
        rom_memory[20203] = 3'b111;
        rom_memory[20204] = 3'b111;
        rom_memory[20205] = 3'b111;
        rom_memory[20206] = 3'b110;
        rom_memory[20207] = 3'b100;
        rom_memory[20208] = 3'b100;
        rom_memory[20209] = 3'b100;
        rom_memory[20210] = 3'b110;
        rom_memory[20211] = 3'b110;
        rom_memory[20212] = 3'b110;
        rom_memory[20213] = 3'b110;
        rom_memory[20214] = 3'b110;
        rom_memory[20215] = 3'b110;
        rom_memory[20216] = 3'b100;
        rom_memory[20217] = 3'b100;
        rom_memory[20218] = 3'b100;
        rom_memory[20219] = 3'b110;
        rom_memory[20220] = 3'b110;
        rom_memory[20221] = 3'b110;
        rom_memory[20222] = 3'b110;
        rom_memory[20223] = 3'b100;
        rom_memory[20224] = 3'b100;
        rom_memory[20225] = 3'b100;
        rom_memory[20226] = 3'b110;
        rom_memory[20227] = 3'b110;
        rom_memory[20228] = 3'b110;
        rom_memory[20229] = 3'b110;
        rom_memory[20230] = 3'b110;
        rom_memory[20231] = 3'b110;
        rom_memory[20232] = 3'b110;
        rom_memory[20233] = 3'b110;
        rom_memory[20234] = 3'b110;
        rom_memory[20235] = 3'b110;
        rom_memory[20236] = 3'b110;
        rom_memory[20237] = 3'b110;
        rom_memory[20238] = 3'b110;
        rom_memory[20239] = 3'b110;
        rom_memory[20240] = 3'b110;
        rom_memory[20241] = 3'b110;
        rom_memory[20242] = 3'b110;
        rom_memory[20243] = 3'b110;
        rom_memory[20244] = 3'b110;
        rom_memory[20245] = 3'b110;
        rom_memory[20246] = 3'b110;
        rom_memory[20247] = 3'b110;
        rom_memory[20248] = 3'b110;
        rom_memory[20249] = 3'b110;
        rom_memory[20250] = 3'b110;
        rom_memory[20251] = 3'b110;
        rom_memory[20252] = 3'b110;
        rom_memory[20253] = 3'b110;
        rom_memory[20254] = 3'b110;
        rom_memory[20255] = 3'b111;
        rom_memory[20256] = 3'b111;
        rom_memory[20257] = 3'b000;
        rom_memory[20258] = 3'b000;
        rom_memory[20259] = 3'b000;
        rom_memory[20260] = 3'b000;
        rom_memory[20261] = 3'b000;
        rom_memory[20262] = 3'b000;
        rom_memory[20263] = 3'b000;
        rom_memory[20264] = 3'b000;
        rom_memory[20265] = 3'b000;
        rom_memory[20266] = 3'b000;
        rom_memory[20267] = 3'b000;
        rom_memory[20268] = 3'b000;
        rom_memory[20269] = 3'b000;
        rom_memory[20270] = 3'b000;
        rom_memory[20271] = 3'b100;
        rom_memory[20272] = 3'b110;
        rom_memory[20273] = 3'b110;
        rom_memory[20274] = 3'b110;
        rom_memory[20275] = 3'b110;
        rom_memory[20276] = 3'b110;
        rom_memory[20277] = 3'b110;
        rom_memory[20278] = 3'b110;
        rom_memory[20279] = 3'b110;
        rom_memory[20280] = 3'b110;
        rom_memory[20281] = 3'b111;
        rom_memory[20282] = 3'b111;
        rom_memory[20283] = 3'b111;
        rom_memory[20284] = 3'b110;
        rom_memory[20285] = 3'b110;
        rom_memory[20286] = 3'b110;
        rom_memory[20287] = 3'b110;
        rom_memory[20288] = 3'b110;
        rom_memory[20289] = 3'b110;
        rom_memory[20290] = 3'b110;
        rom_memory[20291] = 3'b110;
        rom_memory[20292] = 3'b110;
        rom_memory[20293] = 3'b110;
        rom_memory[20294] = 3'b110;
        rom_memory[20295] = 3'b110;
        rom_memory[20296] = 3'b110;
        rom_memory[20297] = 3'b110;
        rom_memory[20298] = 3'b110;
        rom_memory[20299] = 3'b110;
        rom_memory[20300] = 3'b110;
        rom_memory[20301] = 3'b110;
        rom_memory[20302] = 3'b110;
        rom_memory[20303] = 3'b111;
        rom_memory[20304] = 3'b111;
        rom_memory[20305] = 3'b111;
        rom_memory[20306] = 3'b111;
        rom_memory[20307] = 3'b111;
        rom_memory[20308] = 3'b111;
        rom_memory[20309] = 3'b111;
        rom_memory[20310] = 3'b111;
        rom_memory[20311] = 3'b111;
        rom_memory[20312] = 3'b111;
        rom_memory[20313] = 3'b111;
        rom_memory[20314] = 3'b111;
        rom_memory[20315] = 3'b111;
        rom_memory[20316] = 3'b111;
        rom_memory[20317] = 3'b111;
        rom_memory[20318] = 3'b111;
        rom_memory[20319] = 3'b111;
        rom_memory[20320] = 3'b111;
        rom_memory[20321] = 3'b111;
        rom_memory[20322] = 3'b111;
        rom_memory[20323] = 3'b111;
        rom_memory[20324] = 3'b111;
        rom_memory[20325] = 3'b111;
        rom_memory[20326] = 3'b111;
        rom_memory[20327] = 3'b111;
        rom_memory[20328] = 3'b111;
        rom_memory[20329] = 3'b111;
        rom_memory[20330] = 3'b111;
        rom_memory[20331] = 3'b111;
        rom_memory[20332] = 3'b111;
        rom_memory[20333] = 3'b111;
        rom_memory[20334] = 3'b111;
        rom_memory[20335] = 3'b111;
        rom_memory[20336] = 3'b111;
        rom_memory[20337] = 3'b111;
        rom_memory[20338] = 3'b111;
        rom_memory[20339] = 3'b111;
        rom_memory[20340] = 3'b111;
        rom_memory[20341] = 3'b111;
        rom_memory[20342] = 3'b111;
        rom_memory[20343] = 3'b111;
        rom_memory[20344] = 3'b111;
        rom_memory[20345] = 3'b111;
        rom_memory[20346] = 3'b111;
        rom_memory[20347] = 3'b111;
        rom_memory[20348] = 3'b111;
        rom_memory[20349] = 3'b110;
        rom_memory[20350] = 3'b110;
        rom_memory[20351] = 3'b110;
        rom_memory[20352] = 3'b110;
        rom_memory[20353] = 3'b111;
        rom_memory[20354] = 3'b110;
        rom_memory[20355] = 3'b111;
        rom_memory[20356] = 3'b111;
        rom_memory[20357] = 3'b110;
        rom_memory[20358] = 3'b110;
        rom_memory[20359] = 3'b110;
        rom_memory[20360] = 3'b110;
        rom_memory[20361] = 3'b110;
        rom_memory[20362] = 3'b110;
        rom_memory[20363] = 3'b110;
        rom_memory[20364] = 3'b110;
        rom_memory[20365] = 3'b110;
        rom_memory[20366] = 3'b110;
        rom_memory[20367] = 3'b110;
        rom_memory[20368] = 3'b110;
        rom_memory[20369] = 3'b110;
        rom_memory[20370] = 3'b110;
        rom_memory[20371] = 3'b110;
        rom_memory[20372] = 3'b110;
        rom_memory[20373] = 3'b110;
        rom_memory[20374] = 3'b110;
        rom_memory[20375] = 3'b110;
        rom_memory[20376] = 3'b110;
        rom_memory[20377] = 3'b110;
        rom_memory[20378] = 3'b110;
        rom_memory[20379] = 3'b110;
        rom_memory[20380] = 3'b110;
        rom_memory[20381] = 3'b110;
        rom_memory[20382] = 3'b110;
        rom_memory[20383] = 3'b110;
        rom_memory[20384] = 3'b110;
        rom_memory[20385] = 3'b110;
        rom_memory[20386] = 3'b110;
        rom_memory[20387] = 3'b110;
        rom_memory[20388] = 3'b110;
        rom_memory[20389] = 3'b110;
        rom_memory[20390] = 3'b110;
        rom_memory[20391] = 3'b110;
        rom_memory[20392] = 3'b110;
        rom_memory[20393] = 3'b110;
        rom_memory[20394] = 3'b110;
        rom_memory[20395] = 3'b110;
        rom_memory[20396] = 3'b110;
        rom_memory[20397] = 3'b110;
        rom_memory[20398] = 3'b110;
        rom_memory[20399] = 3'b110;
        rom_memory[20400] = 3'b110;
        rom_memory[20401] = 3'b110;
        rom_memory[20402] = 3'b110;
        rom_memory[20403] = 3'b110;
        rom_memory[20404] = 3'b110;
        rom_memory[20405] = 3'b110;
        rom_memory[20406] = 3'b110;
        rom_memory[20407] = 3'b110;
        rom_memory[20408] = 3'b110;
        rom_memory[20409] = 3'b110;
        rom_memory[20410] = 3'b110;
        rom_memory[20411] = 3'b110;
        rom_memory[20412] = 3'b110;
        rom_memory[20413] = 3'b110;
        rom_memory[20414] = 3'b110;
        rom_memory[20415] = 3'b110;
        rom_memory[20416] = 3'b110;
        rom_memory[20417] = 3'b110;
        rom_memory[20418] = 3'b110;
        rom_memory[20419] = 3'b110;
        rom_memory[20420] = 3'b110;
        rom_memory[20421] = 3'b110;
        rom_memory[20422] = 3'b110;
        rom_memory[20423] = 3'b110;
        rom_memory[20424] = 3'b110;
        rom_memory[20425] = 3'b110;
        rom_memory[20426] = 3'b110;
        rom_memory[20427] = 3'b110;
        rom_memory[20428] = 3'b110;
        rom_memory[20429] = 3'b110;
        rom_memory[20430] = 3'b111;
        rom_memory[20431] = 3'b111;
        rom_memory[20432] = 3'b111;
        rom_memory[20433] = 3'b111;
        rom_memory[20434] = 3'b111;
        rom_memory[20435] = 3'b111;
        rom_memory[20436] = 3'b111;
        rom_memory[20437] = 3'b111;
        rom_memory[20438] = 3'b111;
        rom_memory[20439] = 3'b111;
        rom_memory[20440] = 3'b111;
        rom_memory[20441] = 3'b111;
        rom_memory[20442] = 3'b111;
        rom_memory[20443] = 3'b111;
        rom_memory[20444] = 3'b111;
        rom_memory[20445] = 3'b111;
        rom_memory[20446] = 3'b110;
        rom_memory[20447] = 3'b100;
        rom_memory[20448] = 3'b100;
        rom_memory[20449] = 3'b100;
        rom_memory[20450] = 3'b100;
        rom_memory[20451] = 3'b110;
        rom_memory[20452] = 3'b110;
        rom_memory[20453] = 3'b110;
        rom_memory[20454] = 3'b110;
        rom_memory[20455] = 3'b110;
        rom_memory[20456] = 3'b100;
        rom_memory[20457] = 3'b100;
        rom_memory[20458] = 3'b100;
        rom_memory[20459] = 3'b110;
        rom_memory[20460] = 3'b110;
        rom_memory[20461] = 3'b110;
        rom_memory[20462] = 3'b110;
        rom_memory[20463] = 3'b100;
        rom_memory[20464] = 3'b100;
        rom_memory[20465] = 3'b110;
        rom_memory[20466] = 3'b110;
        rom_memory[20467] = 3'b110;
        rom_memory[20468] = 3'b110;
        rom_memory[20469] = 3'b110;
        rom_memory[20470] = 3'b110;
        rom_memory[20471] = 3'b110;
        rom_memory[20472] = 3'b110;
        rom_memory[20473] = 3'b110;
        rom_memory[20474] = 3'b110;
        rom_memory[20475] = 3'b110;
        rom_memory[20476] = 3'b110;
        rom_memory[20477] = 3'b110;
        rom_memory[20478] = 3'b110;
        rom_memory[20479] = 3'b110;
        rom_memory[20480] = 3'b110;
        rom_memory[20481] = 3'b110;
        rom_memory[20482] = 3'b110;
        rom_memory[20483] = 3'b110;
        rom_memory[20484] = 3'b110;
        rom_memory[20485] = 3'b110;
        rom_memory[20486] = 3'b110;
        rom_memory[20487] = 3'b110;
        rom_memory[20488] = 3'b110;
        rom_memory[20489] = 3'b110;
        rom_memory[20490] = 3'b110;
        rom_memory[20491] = 3'b110;
        rom_memory[20492] = 3'b110;
        rom_memory[20493] = 3'b110;
        rom_memory[20494] = 3'b110;
        rom_memory[20495] = 3'b111;
        rom_memory[20496] = 3'b111;
        rom_memory[20497] = 3'b111;
        rom_memory[20498] = 3'b000;
        rom_memory[20499] = 3'b000;
        rom_memory[20500] = 3'b000;
        rom_memory[20501] = 3'b000;
        rom_memory[20502] = 3'b000;
        rom_memory[20503] = 3'b000;
        rom_memory[20504] = 3'b000;
        rom_memory[20505] = 3'b000;
        rom_memory[20506] = 3'b000;
        rom_memory[20507] = 3'b000;
        rom_memory[20508] = 3'b000;
        rom_memory[20509] = 3'b000;
        rom_memory[20510] = 3'b000;
        rom_memory[20511] = 3'b000;
        rom_memory[20512] = 3'b110;
        rom_memory[20513] = 3'b110;
        rom_memory[20514] = 3'b110;
        rom_memory[20515] = 3'b110;
        rom_memory[20516] = 3'b110;
        rom_memory[20517] = 3'b110;
        rom_memory[20518] = 3'b110;
        rom_memory[20519] = 3'b110;
        rom_memory[20520] = 3'b110;
        rom_memory[20521] = 3'b110;
        rom_memory[20522] = 3'b111;
        rom_memory[20523] = 3'b111;
        rom_memory[20524] = 3'b110;
        rom_memory[20525] = 3'b110;
        rom_memory[20526] = 3'b110;
        rom_memory[20527] = 3'b110;
        rom_memory[20528] = 3'b110;
        rom_memory[20529] = 3'b110;
        rom_memory[20530] = 3'b110;
        rom_memory[20531] = 3'b110;
        rom_memory[20532] = 3'b110;
        rom_memory[20533] = 3'b110;
        rom_memory[20534] = 3'b110;
        rom_memory[20535] = 3'b110;
        rom_memory[20536] = 3'b110;
        rom_memory[20537] = 3'b110;
        rom_memory[20538] = 3'b110;
        rom_memory[20539] = 3'b110;
        rom_memory[20540] = 3'b110;
        rom_memory[20541] = 3'b110;
        rom_memory[20542] = 3'b110;
        rom_memory[20543] = 3'b111;
        rom_memory[20544] = 3'b111;
        rom_memory[20545] = 3'b110;
        rom_memory[20546] = 3'b111;
        rom_memory[20547] = 3'b111;
        rom_memory[20548] = 3'b111;
        rom_memory[20549] = 3'b111;
        rom_memory[20550] = 3'b111;
        rom_memory[20551] = 3'b111;
        rom_memory[20552] = 3'b111;
        rom_memory[20553] = 3'b111;
        rom_memory[20554] = 3'b111;
        rom_memory[20555] = 3'b111;
        rom_memory[20556] = 3'b111;
        rom_memory[20557] = 3'b111;
        rom_memory[20558] = 3'b111;
        rom_memory[20559] = 3'b111;
        rom_memory[20560] = 3'b111;
        rom_memory[20561] = 3'b111;
        rom_memory[20562] = 3'b111;
        rom_memory[20563] = 3'b111;
        rom_memory[20564] = 3'b111;
        rom_memory[20565] = 3'b111;
        rom_memory[20566] = 3'b111;
        rom_memory[20567] = 3'b111;
        rom_memory[20568] = 3'b111;
        rom_memory[20569] = 3'b111;
        rom_memory[20570] = 3'b111;
        rom_memory[20571] = 3'b111;
        rom_memory[20572] = 3'b111;
        rom_memory[20573] = 3'b111;
        rom_memory[20574] = 3'b111;
        rom_memory[20575] = 3'b111;
        rom_memory[20576] = 3'b111;
        rom_memory[20577] = 3'b111;
        rom_memory[20578] = 3'b111;
        rom_memory[20579] = 3'b111;
        rom_memory[20580] = 3'b111;
        rom_memory[20581] = 3'b111;
        rom_memory[20582] = 3'b111;
        rom_memory[20583] = 3'b111;
        rom_memory[20584] = 3'b111;
        rom_memory[20585] = 3'b111;
        rom_memory[20586] = 3'b111;
        rom_memory[20587] = 3'b111;
        rom_memory[20588] = 3'b111;
        rom_memory[20589] = 3'b110;
        rom_memory[20590] = 3'b110;
        rom_memory[20591] = 3'b110;
        rom_memory[20592] = 3'b110;
        rom_memory[20593] = 3'b110;
        rom_memory[20594] = 3'b110;
        rom_memory[20595] = 3'b110;
        rom_memory[20596] = 3'b111;
        rom_memory[20597] = 3'b110;
        rom_memory[20598] = 3'b110;
        rom_memory[20599] = 3'b110;
        rom_memory[20600] = 3'b110;
        rom_memory[20601] = 3'b110;
        rom_memory[20602] = 3'b110;
        rom_memory[20603] = 3'b110;
        rom_memory[20604] = 3'b110;
        rom_memory[20605] = 3'b110;
        rom_memory[20606] = 3'b110;
        rom_memory[20607] = 3'b110;
        rom_memory[20608] = 3'b110;
        rom_memory[20609] = 3'b110;
        rom_memory[20610] = 3'b110;
        rom_memory[20611] = 3'b110;
        rom_memory[20612] = 3'b110;
        rom_memory[20613] = 3'b110;
        rom_memory[20614] = 3'b110;
        rom_memory[20615] = 3'b110;
        rom_memory[20616] = 3'b110;
        rom_memory[20617] = 3'b110;
        rom_memory[20618] = 3'b110;
        rom_memory[20619] = 3'b110;
        rom_memory[20620] = 3'b110;
        rom_memory[20621] = 3'b110;
        rom_memory[20622] = 3'b110;
        rom_memory[20623] = 3'b110;
        rom_memory[20624] = 3'b110;
        rom_memory[20625] = 3'b110;
        rom_memory[20626] = 3'b110;
        rom_memory[20627] = 3'b110;
        rom_memory[20628] = 3'b110;
        rom_memory[20629] = 3'b110;
        rom_memory[20630] = 3'b110;
        rom_memory[20631] = 3'b110;
        rom_memory[20632] = 3'b110;
        rom_memory[20633] = 3'b110;
        rom_memory[20634] = 3'b110;
        rom_memory[20635] = 3'b110;
        rom_memory[20636] = 3'b110;
        rom_memory[20637] = 3'b110;
        rom_memory[20638] = 3'b110;
        rom_memory[20639] = 3'b110;
        rom_memory[20640] = 3'b110;
        rom_memory[20641] = 3'b110;
        rom_memory[20642] = 3'b110;
        rom_memory[20643] = 3'b110;
        rom_memory[20644] = 3'b110;
        rom_memory[20645] = 3'b110;
        rom_memory[20646] = 3'b110;
        rom_memory[20647] = 3'b110;
        rom_memory[20648] = 3'b110;
        rom_memory[20649] = 3'b110;
        rom_memory[20650] = 3'b110;
        rom_memory[20651] = 3'b110;
        rom_memory[20652] = 3'b110;
        rom_memory[20653] = 3'b110;
        rom_memory[20654] = 3'b110;
        rom_memory[20655] = 3'b110;
        rom_memory[20656] = 3'b110;
        rom_memory[20657] = 3'b110;
        rom_memory[20658] = 3'b110;
        rom_memory[20659] = 3'b110;
        rom_memory[20660] = 3'b110;
        rom_memory[20661] = 3'b110;
        rom_memory[20662] = 3'b110;
        rom_memory[20663] = 3'b110;
        rom_memory[20664] = 3'b110;
        rom_memory[20665] = 3'b110;
        rom_memory[20666] = 3'b110;
        rom_memory[20667] = 3'b110;
        rom_memory[20668] = 3'b110;
        rom_memory[20669] = 3'b110;
        rom_memory[20670] = 3'b111;
        rom_memory[20671] = 3'b111;
        rom_memory[20672] = 3'b111;
        rom_memory[20673] = 3'b111;
        rom_memory[20674] = 3'b111;
        rom_memory[20675] = 3'b111;
        rom_memory[20676] = 3'b111;
        rom_memory[20677] = 3'b111;
        rom_memory[20678] = 3'b111;
        rom_memory[20679] = 3'b111;
        rom_memory[20680] = 3'b111;
        rom_memory[20681] = 3'b111;
        rom_memory[20682] = 3'b111;
        rom_memory[20683] = 3'b111;
        rom_memory[20684] = 3'b111;
        rom_memory[20685] = 3'b111;
        rom_memory[20686] = 3'b111;
        rom_memory[20687] = 3'b110;
        rom_memory[20688] = 3'b100;
        rom_memory[20689] = 3'b100;
        rom_memory[20690] = 3'b100;
        rom_memory[20691] = 3'b110;
        rom_memory[20692] = 3'b110;
        rom_memory[20693] = 3'b110;
        rom_memory[20694] = 3'b110;
        rom_memory[20695] = 3'b110;
        rom_memory[20696] = 3'b110;
        rom_memory[20697] = 3'b100;
        rom_memory[20698] = 3'b110;
        rom_memory[20699] = 3'b100;
        rom_memory[20700] = 3'b110;
        rom_memory[20701] = 3'b110;
        rom_memory[20702] = 3'b110;
        rom_memory[20703] = 3'b100;
        rom_memory[20704] = 3'b100;
        rom_memory[20705] = 3'b110;
        rom_memory[20706] = 3'b110;
        rom_memory[20707] = 3'b110;
        rom_memory[20708] = 3'b110;
        rom_memory[20709] = 3'b110;
        rom_memory[20710] = 3'b110;
        rom_memory[20711] = 3'b110;
        rom_memory[20712] = 3'b110;
        rom_memory[20713] = 3'b110;
        rom_memory[20714] = 3'b110;
        rom_memory[20715] = 3'b110;
        rom_memory[20716] = 3'b110;
        rom_memory[20717] = 3'b110;
        rom_memory[20718] = 3'b110;
        rom_memory[20719] = 3'b110;
        rom_memory[20720] = 3'b110;
        rom_memory[20721] = 3'b110;
        rom_memory[20722] = 3'b110;
        rom_memory[20723] = 3'b110;
        rom_memory[20724] = 3'b110;
        rom_memory[20725] = 3'b110;
        rom_memory[20726] = 3'b110;
        rom_memory[20727] = 3'b110;
        rom_memory[20728] = 3'b110;
        rom_memory[20729] = 3'b110;
        rom_memory[20730] = 3'b110;
        rom_memory[20731] = 3'b110;
        rom_memory[20732] = 3'b110;
        rom_memory[20733] = 3'b110;
        rom_memory[20734] = 3'b110;
        rom_memory[20735] = 3'b110;
        rom_memory[20736] = 3'b111;
        rom_memory[20737] = 3'b111;
        rom_memory[20738] = 3'b111;
        rom_memory[20739] = 3'b000;
        rom_memory[20740] = 3'b000;
        rom_memory[20741] = 3'b000;
        rom_memory[20742] = 3'b000;
        rom_memory[20743] = 3'b000;
        rom_memory[20744] = 3'b000;
        rom_memory[20745] = 3'b000;
        rom_memory[20746] = 3'b000;
        rom_memory[20747] = 3'b000;
        rom_memory[20748] = 3'b000;
        rom_memory[20749] = 3'b000;
        rom_memory[20750] = 3'b000;
        rom_memory[20751] = 3'b000;
        rom_memory[20752] = 3'b100;
        rom_memory[20753] = 3'b110;
        rom_memory[20754] = 3'b110;
        rom_memory[20755] = 3'b110;
        rom_memory[20756] = 3'b110;
        rom_memory[20757] = 3'b110;
        rom_memory[20758] = 3'b110;
        rom_memory[20759] = 3'b110;
        rom_memory[20760] = 3'b110;
        rom_memory[20761] = 3'b111;
        rom_memory[20762] = 3'b111;
        rom_memory[20763] = 3'b111;
        rom_memory[20764] = 3'b110;
        rom_memory[20765] = 3'b110;
        rom_memory[20766] = 3'b110;
        rom_memory[20767] = 3'b110;
        rom_memory[20768] = 3'b110;
        rom_memory[20769] = 3'b110;
        rom_memory[20770] = 3'b110;
        rom_memory[20771] = 3'b110;
        rom_memory[20772] = 3'b110;
        rom_memory[20773] = 3'b110;
        rom_memory[20774] = 3'b110;
        rom_memory[20775] = 3'b110;
        rom_memory[20776] = 3'b110;
        rom_memory[20777] = 3'b110;
        rom_memory[20778] = 3'b110;
        rom_memory[20779] = 3'b110;
        rom_memory[20780] = 3'b110;
        rom_memory[20781] = 3'b110;
        rom_memory[20782] = 3'b110;
        rom_memory[20783] = 3'b110;
        rom_memory[20784] = 3'b110;
        rom_memory[20785] = 3'b110;
        rom_memory[20786] = 3'b111;
        rom_memory[20787] = 3'b111;
        rom_memory[20788] = 3'b111;
        rom_memory[20789] = 3'b111;
        rom_memory[20790] = 3'b111;
        rom_memory[20791] = 3'b111;
        rom_memory[20792] = 3'b111;
        rom_memory[20793] = 3'b111;
        rom_memory[20794] = 3'b111;
        rom_memory[20795] = 3'b111;
        rom_memory[20796] = 3'b111;
        rom_memory[20797] = 3'b111;
        rom_memory[20798] = 3'b111;
        rom_memory[20799] = 3'b111;
        rom_memory[20800] = 3'b111;
        rom_memory[20801] = 3'b111;
        rom_memory[20802] = 3'b111;
        rom_memory[20803] = 3'b111;
        rom_memory[20804] = 3'b111;
        rom_memory[20805] = 3'b111;
        rom_memory[20806] = 3'b111;
        rom_memory[20807] = 3'b111;
        rom_memory[20808] = 3'b111;
        rom_memory[20809] = 3'b111;
        rom_memory[20810] = 3'b111;
        rom_memory[20811] = 3'b111;
        rom_memory[20812] = 3'b111;
        rom_memory[20813] = 3'b111;
        rom_memory[20814] = 3'b111;
        rom_memory[20815] = 3'b111;
        rom_memory[20816] = 3'b111;
        rom_memory[20817] = 3'b111;
        rom_memory[20818] = 3'b111;
        rom_memory[20819] = 3'b111;
        rom_memory[20820] = 3'b111;
        rom_memory[20821] = 3'b111;
        rom_memory[20822] = 3'b111;
        rom_memory[20823] = 3'b111;
        rom_memory[20824] = 3'b111;
        rom_memory[20825] = 3'b111;
        rom_memory[20826] = 3'b111;
        rom_memory[20827] = 3'b111;
        rom_memory[20828] = 3'b110;
        rom_memory[20829] = 3'b110;
        rom_memory[20830] = 3'b110;
        rom_memory[20831] = 3'b110;
        rom_memory[20832] = 3'b110;
        rom_memory[20833] = 3'b110;
        rom_memory[20834] = 3'b110;
        rom_memory[20835] = 3'b110;
        rom_memory[20836] = 3'b110;
        rom_memory[20837] = 3'b110;
        rom_memory[20838] = 3'b110;
        rom_memory[20839] = 3'b110;
        rom_memory[20840] = 3'b110;
        rom_memory[20841] = 3'b110;
        rom_memory[20842] = 3'b110;
        rom_memory[20843] = 3'b110;
        rom_memory[20844] = 3'b110;
        rom_memory[20845] = 3'b110;
        rom_memory[20846] = 3'b110;
        rom_memory[20847] = 3'b110;
        rom_memory[20848] = 3'b110;
        rom_memory[20849] = 3'b110;
        rom_memory[20850] = 3'b110;
        rom_memory[20851] = 3'b110;
        rom_memory[20852] = 3'b110;
        rom_memory[20853] = 3'b110;
        rom_memory[20854] = 3'b110;
        rom_memory[20855] = 3'b110;
        rom_memory[20856] = 3'b110;
        rom_memory[20857] = 3'b110;
        rom_memory[20858] = 3'b110;
        rom_memory[20859] = 3'b110;
        rom_memory[20860] = 3'b110;
        rom_memory[20861] = 3'b110;
        rom_memory[20862] = 3'b110;
        rom_memory[20863] = 3'b110;
        rom_memory[20864] = 3'b110;
        rom_memory[20865] = 3'b110;
        rom_memory[20866] = 3'b110;
        rom_memory[20867] = 3'b110;
        rom_memory[20868] = 3'b110;
        rom_memory[20869] = 3'b110;
        rom_memory[20870] = 3'b110;
        rom_memory[20871] = 3'b110;
        rom_memory[20872] = 3'b110;
        rom_memory[20873] = 3'b110;
        rom_memory[20874] = 3'b110;
        rom_memory[20875] = 3'b110;
        rom_memory[20876] = 3'b110;
        rom_memory[20877] = 3'b110;
        rom_memory[20878] = 3'b110;
        rom_memory[20879] = 3'b110;
        rom_memory[20880] = 3'b110;
        rom_memory[20881] = 3'b110;
        rom_memory[20882] = 3'b110;
        rom_memory[20883] = 3'b110;
        rom_memory[20884] = 3'b110;
        rom_memory[20885] = 3'b110;
        rom_memory[20886] = 3'b110;
        rom_memory[20887] = 3'b110;
        rom_memory[20888] = 3'b110;
        rom_memory[20889] = 3'b110;
        rom_memory[20890] = 3'b110;
        rom_memory[20891] = 3'b110;
        rom_memory[20892] = 3'b110;
        rom_memory[20893] = 3'b110;
        rom_memory[20894] = 3'b110;
        rom_memory[20895] = 3'b110;
        rom_memory[20896] = 3'b110;
        rom_memory[20897] = 3'b110;
        rom_memory[20898] = 3'b110;
        rom_memory[20899] = 3'b110;
        rom_memory[20900] = 3'b110;
        rom_memory[20901] = 3'b110;
        rom_memory[20902] = 3'b110;
        rom_memory[20903] = 3'b110;
        rom_memory[20904] = 3'b110;
        rom_memory[20905] = 3'b110;
        rom_memory[20906] = 3'b110;
        rom_memory[20907] = 3'b110;
        rom_memory[20908] = 3'b110;
        rom_memory[20909] = 3'b110;
        rom_memory[20910] = 3'b111;
        rom_memory[20911] = 3'b111;
        rom_memory[20912] = 3'b111;
        rom_memory[20913] = 3'b111;
        rom_memory[20914] = 3'b111;
        rom_memory[20915] = 3'b111;
        rom_memory[20916] = 3'b111;
        rom_memory[20917] = 3'b111;
        rom_memory[20918] = 3'b111;
        rom_memory[20919] = 3'b111;
        rom_memory[20920] = 3'b111;
        rom_memory[20921] = 3'b111;
        rom_memory[20922] = 3'b111;
        rom_memory[20923] = 3'b111;
        rom_memory[20924] = 3'b111;
        rom_memory[20925] = 3'b111;
        rom_memory[20926] = 3'b111;
        rom_memory[20927] = 3'b110;
        rom_memory[20928] = 3'b100;
        rom_memory[20929] = 3'b100;
        rom_memory[20930] = 3'b100;
        rom_memory[20931] = 3'b110;
        rom_memory[20932] = 3'b110;
        rom_memory[20933] = 3'b110;
        rom_memory[20934] = 3'b110;
        rom_memory[20935] = 3'b110;
        rom_memory[20936] = 3'b110;
        rom_memory[20937] = 3'b110;
        rom_memory[20938] = 3'b100;
        rom_memory[20939] = 3'b100;
        rom_memory[20940] = 3'b110;
        rom_memory[20941] = 3'b110;
        rom_memory[20942] = 3'b110;
        rom_memory[20943] = 3'b110;
        rom_memory[20944] = 3'b100;
        rom_memory[20945] = 3'b110;
        rom_memory[20946] = 3'b100;
        rom_memory[20947] = 3'b110;
        rom_memory[20948] = 3'b110;
        rom_memory[20949] = 3'b110;
        rom_memory[20950] = 3'b110;
        rom_memory[20951] = 3'b110;
        rom_memory[20952] = 3'b110;
        rom_memory[20953] = 3'b110;
        rom_memory[20954] = 3'b110;
        rom_memory[20955] = 3'b110;
        rom_memory[20956] = 3'b110;
        rom_memory[20957] = 3'b110;
        rom_memory[20958] = 3'b110;
        rom_memory[20959] = 3'b110;
        rom_memory[20960] = 3'b110;
        rom_memory[20961] = 3'b110;
        rom_memory[20962] = 3'b110;
        rom_memory[20963] = 3'b110;
        rom_memory[20964] = 3'b110;
        rom_memory[20965] = 3'b110;
        rom_memory[20966] = 3'b110;
        rom_memory[20967] = 3'b110;
        rom_memory[20968] = 3'b110;
        rom_memory[20969] = 3'b110;
        rom_memory[20970] = 3'b110;
        rom_memory[20971] = 3'b110;
        rom_memory[20972] = 3'b110;
        rom_memory[20973] = 3'b110;
        rom_memory[20974] = 3'b110;
        rom_memory[20975] = 3'b110;
        rom_memory[20976] = 3'b111;
        rom_memory[20977] = 3'b111;
        rom_memory[20978] = 3'b111;
        rom_memory[20979] = 3'b111;
        rom_memory[20980] = 3'b110;
        rom_memory[20981] = 3'b000;
        rom_memory[20982] = 3'b000;
        rom_memory[20983] = 3'b000;
        rom_memory[20984] = 3'b000;
        rom_memory[20985] = 3'b000;
        rom_memory[20986] = 3'b000;
        rom_memory[20987] = 3'b000;
        rom_memory[20988] = 3'b000;
        rom_memory[20989] = 3'b000;
        rom_memory[20990] = 3'b000;
        rom_memory[20991] = 3'b000;
        rom_memory[20992] = 3'b000;
        rom_memory[20993] = 3'b110;
        rom_memory[20994] = 3'b100;
        rom_memory[20995] = 3'b110;
        rom_memory[20996] = 3'b110;
        rom_memory[20997] = 3'b110;
        rom_memory[20998] = 3'b110;
        rom_memory[20999] = 3'b110;
        rom_memory[21000] = 3'b110;
        rom_memory[21001] = 3'b110;
        rom_memory[21002] = 3'b111;
        rom_memory[21003] = 3'b111;
        rom_memory[21004] = 3'b111;
        rom_memory[21005] = 3'b110;
        rom_memory[21006] = 3'b110;
        rom_memory[21007] = 3'b110;
        rom_memory[21008] = 3'b110;
        rom_memory[21009] = 3'b110;
        rom_memory[21010] = 3'b110;
        rom_memory[21011] = 3'b110;
        rom_memory[21012] = 3'b110;
        rom_memory[21013] = 3'b110;
        rom_memory[21014] = 3'b110;
        rom_memory[21015] = 3'b110;
        rom_memory[21016] = 3'b110;
        rom_memory[21017] = 3'b110;
        rom_memory[21018] = 3'b110;
        rom_memory[21019] = 3'b110;
        rom_memory[21020] = 3'b110;
        rom_memory[21021] = 3'b110;
        rom_memory[21022] = 3'b110;
        rom_memory[21023] = 3'b110;
        rom_memory[21024] = 3'b110;
        rom_memory[21025] = 3'b110;
        rom_memory[21026] = 3'b110;
        rom_memory[21027] = 3'b111;
        rom_memory[21028] = 3'b111;
        rom_memory[21029] = 3'b111;
        rom_memory[21030] = 3'b111;
        rom_memory[21031] = 3'b111;
        rom_memory[21032] = 3'b111;
        rom_memory[21033] = 3'b111;
        rom_memory[21034] = 3'b111;
        rom_memory[21035] = 3'b111;
        rom_memory[21036] = 3'b111;
        rom_memory[21037] = 3'b111;
        rom_memory[21038] = 3'b111;
        rom_memory[21039] = 3'b111;
        rom_memory[21040] = 3'b111;
        rom_memory[21041] = 3'b111;
        rom_memory[21042] = 3'b111;
        rom_memory[21043] = 3'b111;
        rom_memory[21044] = 3'b111;
        rom_memory[21045] = 3'b111;
        rom_memory[21046] = 3'b111;
        rom_memory[21047] = 3'b111;
        rom_memory[21048] = 3'b111;
        rom_memory[21049] = 3'b111;
        rom_memory[21050] = 3'b111;
        rom_memory[21051] = 3'b111;
        rom_memory[21052] = 3'b111;
        rom_memory[21053] = 3'b111;
        rom_memory[21054] = 3'b111;
        rom_memory[21055] = 3'b111;
        rom_memory[21056] = 3'b111;
        rom_memory[21057] = 3'b111;
        rom_memory[21058] = 3'b111;
        rom_memory[21059] = 3'b111;
        rom_memory[21060] = 3'b111;
        rom_memory[21061] = 3'b111;
        rom_memory[21062] = 3'b111;
        rom_memory[21063] = 3'b111;
        rom_memory[21064] = 3'b111;
        rom_memory[21065] = 3'b111;
        rom_memory[21066] = 3'b111;
        rom_memory[21067] = 3'b111;
        rom_memory[21068] = 3'b111;
        rom_memory[21069] = 3'b111;
        rom_memory[21070] = 3'b110;
        rom_memory[21071] = 3'b110;
        rom_memory[21072] = 3'b110;
        rom_memory[21073] = 3'b110;
        rom_memory[21074] = 3'b110;
        rom_memory[21075] = 3'b110;
        rom_memory[21076] = 3'b110;
        rom_memory[21077] = 3'b110;
        rom_memory[21078] = 3'b110;
        rom_memory[21079] = 3'b110;
        rom_memory[21080] = 3'b110;
        rom_memory[21081] = 3'b110;
        rom_memory[21082] = 3'b110;
        rom_memory[21083] = 3'b110;
        rom_memory[21084] = 3'b110;
        rom_memory[21085] = 3'b110;
        rom_memory[21086] = 3'b110;
        rom_memory[21087] = 3'b110;
        rom_memory[21088] = 3'b110;
        rom_memory[21089] = 3'b110;
        rom_memory[21090] = 3'b110;
        rom_memory[21091] = 3'b110;
        rom_memory[21092] = 3'b110;
        rom_memory[21093] = 3'b110;
        rom_memory[21094] = 3'b110;
        rom_memory[21095] = 3'b110;
        rom_memory[21096] = 3'b110;
        rom_memory[21097] = 3'b110;
        rom_memory[21098] = 3'b110;
        rom_memory[21099] = 3'b110;
        rom_memory[21100] = 3'b110;
        rom_memory[21101] = 3'b110;
        rom_memory[21102] = 3'b110;
        rom_memory[21103] = 3'b110;
        rom_memory[21104] = 3'b110;
        rom_memory[21105] = 3'b110;
        rom_memory[21106] = 3'b110;
        rom_memory[21107] = 3'b110;
        rom_memory[21108] = 3'b110;
        rom_memory[21109] = 3'b110;
        rom_memory[21110] = 3'b110;
        rom_memory[21111] = 3'b110;
        rom_memory[21112] = 3'b110;
        rom_memory[21113] = 3'b110;
        rom_memory[21114] = 3'b110;
        rom_memory[21115] = 3'b110;
        rom_memory[21116] = 3'b110;
        rom_memory[21117] = 3'b110;
        rom_memory[21118] = 3'b110;
        rom_memory[21119] = 3'b110;
        rom_memory[21120] = 3'b110;
        rom_memory[21121] = 3'b110;
        rom_memory[21122] = 3'b110;
        rom_memory[21123] = 3'b110;
        rom_memory[21124] = 3'b110;
        rom_memory[21125] = 3'b110;
        rom_memory[21126] = 3'b110;
        rom_memory[21127] = 3'b110;
        rom_memory[21128] = 3'b110;
        rom_memory[21129] = 3'b110;
        rom_memory[21130] = 3'b110;
        rom_memory[21131] = 3'b110;
        rom_memory[21132] = 3'b110;
        rom_memory[21133] = 3'b110;
        rom_memory[21134] = 3'b110;
        rom_memory[21135] = 3'b110;
        rom_memory[21136] = 3'b110;
        rom_memory[21137] = 3'b110;
        rom_memory[21138] = 3'b110;
        rom_memory[21139] = 3'b110;
        rom_memory[21140] = 3'b110;
        rom_memory[21141] = 3'b110;
        rom_memory[21142] = 3'b110;
        rom_memory[21143] = 3'b110;
        rom_memory[21144] = 3'b110;
        rom_memory[21145] = 3'b110;
        rom_memory[21146] = 3'b110;
        rom_memory[21147] = 3'b110;
        rom_memory[21148] = 3'b110;
        rom_memory[21149] = 3'b110;
        rom_memory[21150] = 3'b110;
        rom_memory[21151] = 3'b111;
        rom_memory[21152] = 3'b111;
        rom_memory[21153] = 3'b111;
        rom_memory[21154] = 3'b111;
        rom_memory[21155] = 3'b111;
        rom_memory[21156] = 3'b111;
        rom_memory[21157] = 3'b111;
        rom_memory[21158] = 3'b111;
        rom_memory[21159] = 3'b111;
        rom_memory[21160] = 3'b111;
        rom_memory[21161] = 3'b111;
        rom_memory[21162] = 3'b111;
        rom_memory[21163] = 3'b111;
        rom_memory[21164] = 3'b111;
        rom_memory[21165] = 3'b111;
        rom_memory[21166] = 3'b111;
        rom_memory[21167] = 3'b110;
        rom_memory[21168] = 3'b100;
        rom_memory[21169] = 3'b100;
        rom_memory[21170] = 3'b100;
        rom_memory[21171] = 3'b110;
        rom_memory[21172] = 3'b110;
        rom_memory[21173] = 3'b110;
        rom_memory[21174] = 3'b110;
        rom_memory[21175] = 3'b110;
        rom_memory[21176] = 3'b100;
        rom_memory[21177] = 3'b110;
        rom_memory[21178] = 3'b100;
        rom_memory[21179] = 3'b100;
        rom_memory[21180] = 3'b110;
        rom_memory[21181] = 3'b110;
        rom_memory[21182] = 3'b110;
        rom_memory[21183] = 3'b110;
        rom_memory[21184] = 3'b100;
        rom_memory[21185] = 3'b100;
        rom_memory[21186] = 3'b110;
        rom_memory[21187] = 3'b110;
        rom_memory[21188] = 3'b110;
        rom_memory[21189] = 3'b100;
        rom_memory[21190] = 3'b110;
        rom_memory[21191] = 3'b110;
        rom_memory[21192] = 3'b110;
        rom_memory[21193] = 3'b110;
        rom_memory[21194] = 3'b110;
        rom_memory[21195] = 3'b110;
        rom_memory[21196] = 3'b110;
        rom_memory[21197] = 3'b110;
        rom_memory[21198] = 3'b110;
        rom_memory[21199] = 3'b110;
        rom_memory[21200] = 3'b110;
        rom_memory[21201] = 3'b110;
        rom_memory[21202] = 3'b110;
        rom_memory[21203] = 3'b110;
        rom_memory[21204] = 3'b110;
        rom_memory[21205] = 3'b110;
        rom_memory[21206] = 3'b110;
        rom_memory[21207] = 3'b110;
        rom_memory[21208] = 3'b110;
        rom_memory[21209] = 3'b110;
        rom_memory[21210] = 3'b110;
        rom_memory[21211] = 3'b110;
        rom_memory[21212] = 3'b110;
        rom_memory[21213] = 3'b110;
        rom_memory[21214] = 3'b110;
        rom_memory[21215] = 3'b110;
        rom_memory[21216] = 3'b110;
        rom_memory[21217] = 3'b111;
        rom_memory[21218] = 3'b111;
        rom_memory[21219] = 3'b111;
        rom_memory[21220] = 3'b111;
        rom_memory[21221] = 3'b111;
        rom_memory[21222] = 3'b100;
        rom_memory[21223] = 3'b000;
        rom_memory[21224] = 3'b000;
        rom_memory[21225] = 3'b000;
        rom_memory[21226] = 3'b000;
        rom_memory[21227] = 3'b000;
        rom_memory[21228] = 3'b000;
        rom_memory[21229] = 3'b000;
        rom_memory[21230] = 3'b000;
        rom_memory[21231] = 3'b000;
        rom_memory[21232] = 3'b000;
        rom_memory[21233] = 3'b000;
        rom_memory[21234] = 3'b110;
        rom_memory[21235] = 3'b100;
        rom_memory[21236] = 3'b110;
        rom_memory[21237] = 3'b110;
        rom_memory[21238] = 3'b110;
        rom_memory[21239] = 3'b110;
        rom_memory[21240] = 3'b110;
        rom_memory[21241] = 3'b110;
        rom_memory[21242] = 3'b110;
        rom_memory[21243] = 3'b111;
        rom_memory[21244] = 3'b111;
        rom_memory[21245] = 3'b111;
        rom_memory[21246] = 3'b110;
        rom_memory[21247] = 3'b110;
        rom_memory[21248] = 3'b110;
        rom_memory[21249] = 3'b110;
        rom_memory[21250] = 3'b110;
        rom_memory[21251] = 3'b110;
        rom_memory[21252] = 3'b110;
        rom_memory[21253] = 3'b110;
        rom_memory[21254] = 3'b110;
        rom_memory[21255] = 3'b110;
        rom_memory[21256] = 3'b110;
        rom_memory[21257] = 3'b110;
        rom_memory[21258] = 3'b110;
        rom_memory[21259] = 3'b110;
        rom_memory[21260] = 3'b110;
        rom_memory[21261] = 3'b110;
        rom_memory[21262] = 3'b110;
        rom_memory[21263] = 3'b110;
        rom_memory[21264] = 3'b110;
        rom_memory[21265] = 3'b110;
        rom_memory[21266] = 3'b110;
        rom_memory[21267] = 3'b111;
        rom_memory[21268] = 3'b111;
        rom_memory[21269] = 3'b111;
        rom_memory[21270] = 3'b111;
        rom_memory[21271] = 3'b111;
        rom_memory[21272] = 3'b111;
        rom_memory[21273] = 3'b111;
        rom_memory[21274] = 3'b111;
        rom_memory[21275] = 3'b111;
        rom_memory[21276] = 3'b111;
        rom_memory[21277] = 3'b111;
        rom_memory[21278] = 3'b111;
        rom_memory[21279] = 3'b111;
        rom_memory[21280] = 3'b111;
        rom_memory[21281] = 3'b111;
        rom_memory[21282] = 3'b111;
        rom_memory[21283] = 3'b111;
        rom_memory[21284] = 3'b111;
        rom_memory[21285] = 3'b111;
        rom_memory[21286] = 3'b111;
        rom_memory[21287] = 3'b111;
        rom_memory[21288] = 3'b111;
        rom_memory[21289] = 3'b111;
        rom_memory[21290] = 3'b111;
        rom_memory[21291] = 3'b111;
        rom_memory[21292] = 3'b111;
        rom_memory[21293] = 3'b111;
        rom_memory[21294] = 3'b111;
        rom_memory[21295] = 3'b111;
        rom_memory[21296] = 3'b111;
        rom_memory[21297] = 3'b111;
        rom_memory[21298] = 3'b111;
        rom_memory[21299] = 3'b111;
        rom_memory[21300] = 3'b111;
        rom_memory[21301] = 3'b111;
        rom_memory[21302] = 3'b111;
        rom_memory[21303] = 3'b111;
        rom_memory[21304] = 3'b111;
        rom_memory[21305] = 3'b110;
        rom_memory[21306] = 3'b111;
        rom_memory[21307] = 3'b111;
        rom_memory[21308] = 3'b111;
        rom_memory[21309] = 3'b111;
        rom_memory[21310] = 3'b111;
        rom_memory[21311] = 3'b110;
        rom_memory[21312] = 3'b110;
        rom_memory[21313] = 3'b110;
        rom_memory[21314] = 3'b110;
        rom_memory[21315] = 3'b110;
        rom_memory[21316] = 3'b110;
        rom_memory[21317] = 3'b110;
        rom_memory[21318] = 3'b110;
        rom_memory[21319] = 3'b110;
        rom_memory[21320] = 3'b110;
        rom_memory[21321] = 3'b110;
        rom_memory[21322] = 3'b110;
        rom_memory[21323] = 3'b110;
        rom_memory[21324] = 3'b110;
        rom_memory[21325] = 3'b110;
        rom_memory[21326] = 3'b110;
        rom_memory[21327] = 3'b110;
        rom_memory[21328] = 3'b110;
        rom_memory[21329] = 3'b110;
        rom_memory[21330] = 3'b110;
        rom_memory[21331] = 3'b110;
        rom_memory[21332] = 3'b110;
        rom_memory[21333] = 3'b110;
        rom_memory[21334] = 3'b110;
        rom_memory[21335] = 3'b110;
        rom_memory[21336] = 3'b110;
        rom_memory[21337] = 3'b110;
        rom_memory[21338] = 3'b110;
        rom_memory[21339] = 3'b110;
        rom_memory[21340] = 3'b110;
        rom_memory[21341] = 3'b110;
        rom_memory[21342] = 3'b110;
        rom_memory[21343] = 3'b110;
        rom_memory[21344] = 3'b110;
        rom_memory[21345] = 3'b110;
        rom_memory[21346] = 3'b110;
        rom_memory[21347] = 3'b110;
        rom_memory[21348] = 3'b110;
        rom_memory[21349] = 3'b110;
        rom_memory[21350] = 3'b110;
        rom_memory[21351] = 3'b110;
        rom_memory[21352] = 3'b110;
        rom_memory[21353] = 3'b110;
        rom_memory[21354] = 3'b110;
        rom_memory[21355] = 3'b110;
        rom_memory[21356] = 3'b110;
        rom_memory[21357] = 3'b110;
        rom_memory[21358] = 3'b110;
        rom_memory[21359] = 3'b110;
        rom_memory[21360] = 3'b110;
        rom_memory[21361] = 3'b110;
        rom_memory[21362] = 3'b110;
        rom_memory[21363] = 3'b110;
        rom_memory[21364] = 3'b110;
        rom_memory[21365] = 3'b110;
        rom_memory[21366] = 3'b110;
        rom_memory[21367] = 3'b110;
        rom_memory[21368] = 3'b110;
        rom_memory[21369] = 3'b110;
        rom_memory[21370] = 3'b110;
        rom_memory[21371] = 3'b110;
        rom_memory[21372] = 3'b110;
        rom_memory[21373] = 3'b110;
        rom_memory[21374] = 3'b110;
        rom_memory[21375] = 3'b110;
        rom_memory[21376] = 3'b110;
        rom_memory[21377] = 3'b110;
        rom_memory[21378] = 3'b110;
        rom_memory[21379] = 3'b110;
        rom_memory[21380] = 3'b110;
        rom_memory[21381] = 3'b110;
        rom_memory[21382] = 3'b110;
        rom_memory[21383] = 3'b110;
        rom_memory[21384] = 3'b110;
        rom_memory[21385] = 3'b110;
        rom_memory[21386] = 3'b110;
        rom_memory[21387] = 3'b110;
        rom_memory[21388] = 3'b110;
        rom_memory[21389] = 3'b110;
        rom_memory[21390] = 3'b110;
        rom_memory[21391] = 3'b111;
        rom_memory[21392] = 3'b111;
        rom_memory[21393] = 3'b111;
        rom_memory[21394] = 3'b111;
        rom_memory[21395] = 3'b111;
        rom_memory[21396] = 3'b111;
        rom_memory[21397] = 3'b111;
        rom_memory[21398] = 3'b111;
        rom_memory[21399] = 3'b111;
        rom_memory[21400] = 3'b111;
        rom_memory[21401] = 3'b111;
        rom_memory[21402] = 3'b111;
        rom_memory[21403] = 3'b111;
        rom_memory[21404] = 3'b111;
        rom_memory[21405] = 3'b111;
        rom_memory[21406] = 3'b110;
        rom_memory[21407] = 3'b110;
        rom_memory[21408] = 3'b100;
        rom_memory[21409] = 3'b100;
        rom_memory[21410] = 3'b110;
        rom_memory[21411] = 3'b110;
        rom_memory[21412] = 3'b110;
        rom_memory[21413] = 3'b110;
        rom_memory[21414] = 3'b110;
        rom_memory[21415] = 3'b110;
        rom_memory[21416] = 3'b100;
        rom_memory[21417] = 3'b110;
        rom_memory[21418] = 3'b110;
        rom_memory[21419] = 3'b100;
        rom_memory[21420] = 3'b110;
        rom_memory[21421] = 3'b110;
        rom_memory[21422] = 3'b100;
        rom_memory[21423] = 3'b110;
        rom_memory[21424] = 3'b110;
        rom_memory[21425] = 3'b110;
        rom_memory[21426] = 3'b110;
        rom_memory[21427] = 3'b110;
        rom_memory[21428] = 3'b110;
        rom_memory[21429] = 3'b110;
        rom_memory[21430] = 3'b110;
        rom_memory[21431] = 3'b110;
        rom_memory[21432] = 3'b110;
        rom_memory[21433] = 3'b110;
        rom_memory[21434] = 3'b110;
        rom_memory[21435] = 3'b110;
        rom_memory[21436] = 3'b110;
        rom_memory[21437] = 3'b110;
        rom_memory[21438] = 3'b110;
        rom_memory[21439] = 3'b110;
        rom_memory[21440] = 3'b110;
        rom_memory[21441] = 3'b110;
        rom_memory[21442] = 3'b110;
        rom_memory[21443] = 3'b110;
        rom_memory[21444] = 3'b110;
        rom_memory[21445] = 3'b110;
        rom_memory[21446] = 3'b110;
        rom_memory[21447] = 3'b110;
        rom_memory[21448] = 3'b110;
        rom_memory[21449] = 3'b110;
        rom_memory[21450] = 3'b110;
        rom_memory[21451] = 3'b110;
        rom_memory[21452] = 3'b110;
        rom_memory[21453] = 3'b110;
        rom_memory[21454] = 3'b110;
        rom_memory[21455] = 3'b110;
        rom_memory[21456] = 3'b110;
        rom_memory[21457] = 3'b111;
        rom_memory[21458] = 3'b111;
        rom_memory[21459] = 3'b111;
        rom_memory[21460] = 3'b111;
        rom_memory[21461] = 3'b111;
        rom_memory[21462] = 3'b111;
        rom_memory[21463] = 3'b111;
        rom_memory[21464] = 3'b000;
        rom_memory[21465] = 3'b000;
        rom_memory[21466] = 3'b000;
        rom_memory[21467] = 3'b000;
        rom_memory[21468] = 3'b000;
        rom_memory[21469] = 3'b000;
        rom_memory[21470] = 3'b000;
        rom_memory[21471] = 3'b000;
        rom_memory[21472] = 3'b000;
        rom_memory[21473] = 3'b100;
        rom_memory[21474] = 3'b100;
        rom_memory[21475] = 3'b110;
        rom_memory[21476] = 3'b100;
        rom_memory[21477] = 3'b110;
        rom_memory[21478] = 3'b110;
        rom_memory[21479] = 3'b110;
        rom_memory[21480] = 3'b110;
        rom_memory[21481] = 3'b110;
        rom_memory[21482] = 3'b110;
        rom_memory[21483] = 3'b110;
        rom_memory[21484] = 3'b111;
        rom_memory[21485] = 3'b111;
        rom_memory[21486] = 3'b111;
        rom_memory[21487] = 3'b110;
        rom_memory[21488] = 3'b110;
        rom_memory[21489] = 3'b110;
        rom_memory[21490] = 3'b110;
        rom_memory[21491] = 3'b110;
        rom_memory[21492] = 3'b110;
        rom_memory[21493] = 3'b110;
        rom_memory[21494] = 3'b110;
        rom_memory[21495] = 3'b110;
        rom_memory[21496] = 3'b110;
        rom_memory[21497] = 3'b110;
        rom_memory[21498] = 3'b110;
        rom_memory[21499] = 3'b110;
        rom_memory[21500] = 3'b110;
        rom_memory[21501] = 3'b110;
        rom_memory[21502] = 3'b110;
        rom_memory[21503] = 3'b110;
        rom_memory[21504] = 3'b110;
        rom_memory[21505] = 3'b110;
        rom_memory[21506] = 3'b110;
        rom_memory[21507] = 3'b111;
        rom_memory[21508] = 3'b111;
        rom_memory[21509] = 3'b111;
        rom_memory[21510] = 3'b111;
        rom_memory[21511] = 3'b111;
        rom_memory[21512] = 3'b111;
        rom_memory[21513] = 3'b111;
        rom_memory[21514] = 3'b111;
        rom_memory[21515] = 3'b111;
        rom_memory[21516] = 3'b111;
        rom_memory[21517] = 3'b111;
        rom_memory[21518] = 3'b111;
        rom_memory[21519] = 3'b111;
        rom_memory[21520] = 3'b111;
        rom_memory[21521] = 3'b111;
        rom_memory[21522] = 3'b111;
        rom_memory[21523] = 3'b111;
        rom_memory[21524] = 3'b111;
        rom_memory[21525] = 3'b111;
        rom_memory[21526] = 3'b111;
        rom_memory[21527] = 3'b111;
        rom_memory[21528] = 3'b111;
        rom_memory[21529] = 3'b111;
        rom_memory[21530] = 3'b111;
        rom_memory[21531] = 3'b111;
        rom_memory[21532] = 3'b111;
        rom_memory[21533] = 3'b111;
        rom_memory[21534] = 3'b111;
        rom_memory[21535] = 3'b111;
        rom_memory[21536] = 3'b111;
        rom_memory[21537] = 3'b111;
        rom_memory[21538] = 3'b111;
        rom_memory[21539] = 3'b111;
        rom_memory[21540] = 3'b111;
        rom_memory[21541] = 3'b111;
        rom_memory[21542] = 3'b111;
        rom_memory[21543] = 3'b111;
        rom_memory[21544] = 3'b111;
        rom_memory[21545] = 3'b111;
        rom_memory[21546] = 3'b111;
        rom_memory[21547] = 3'b111;
        rom_memory[21548] = 3'b111;
        rom_memory[21549] = 3'b111;
        rom_memory[21550] = 3'b111;
        rom_memory[21551] = 3'b110;
        rom_memory[21552] = 3'b110;
        rom_memory[21553] = 3'b110;
        rom_memory[21554] = 3'b110;
        rom_memory[21555] = 3'b110;
        rom_memory[21556] = 3'b111;
        rom_memory[21557] = 3'b110;
        rom_memory[21558] = 3'b110;
        rom_memory[21559] = 3'b110;
        rom_memory[21560] = 3'b110;
        rom_memory[21561] = 3'b110;
        rom_memory[21562] = 3'b110;
        rom_memory[21563] = 3'b110;
        rom_memory[21564] = 3'b110;
        rom_memory[21565] = 3'b110;
        rom_memory[21566] = 3'b111;
        rom_memory[21567] = 3'b110;
        rom_memory[21568] = 3'b110;
        rom_memory[21569] = 3'b110;
        rom_memory[21570] = 3'b110;
        rom_memory[21571] = 3'b110;
        rom_memory[21572] = 3'b110;
        rom_memory[21573] = 3'b110;
        rom_memory[21574] = 3'b110;
        rom_memory[21575] = 3'b110;
        rom_memory[21576] = 3'b110;
        rom_memory[21577] = 3'b110;
        rom_memory[21578] = 3'b110;
        rom_memory[21579] = 3'b110;
        rom_memory[21580] = 3'b110;
        rom_memory[21581] = 3'b110;
        rom_memory[21582] = 3'b110;
        rom_memory[21583] = 3'b110;
        rom_memory[21584] = 3'b110;
        rom_memory[21585] = 3'b110;
        rom_memory[21586] = 3'b110;
        rom_memory[21587] = 3'b110;
        rom_memory[21588] = 3'b110;
        rom_memory[21589] = 3'b110;
        rom_memory[21590] = 3'b110;
        rom_memory[21591] = 3'b110;
        rom_memory[21592] = 3'b110;
        rom_memory[21593] = 3'b110;
        rom_memory[21594] = 3'b110;
        rom_memory[21595] = 3'b110;
        rom_memory[21596] = 3'b110;
        rom_memory[21597] = 3'b110;
        rom_memory[21598] = 3'b110;
        rom_memory[21599] = 3'b110;
        rom_memory[21600] = 3'b110;
        rom_memory[21601] = 3'b110;
        rom_memory[21602] = 3'b110;
        rom_memory[21603] = 3'b110;
        rom_memory[21604] = 3'b110;
        rom_memory[21605] = 3'b110;
        rom_memory[21606] = 3'b110;
        rom_memory[21607] = 3'b110;
        rom_memory[21608] = 3'b110;
        rom_memory[21609] = 3'b110;
        rom_memory[21610] = 3'b110;
        rom_memory[21611] = 3'b110;
        rom_memory[21612] = 3'b110;
        rom_memory[21613] = 3'b110;
        rom_memory[21614] = 3'b110;
        rom_memory[21615] = 3'b110;
        rom_memory[21616] = 3'b110;
        rom_memory[21617] = 3'b110;
        rom_memory[21618] = 3'b110;
        rom_memory[21619] = 3'b110;
        rom_memory[21620] = 3'b110;
        rom_memory[21621] = 3'b110;
        rom_memory[21622] = 3'b110;
        rom_memory[21623] = 3'b110;
        rom_memory[21624] = 3'b110;
        rom_memory[21625] = 3'b110;
        rom_memory[21626] = 3'b110;
        rom_memory[21627] = 3'b110;
        rom_memory[21628] = 3'b110;
        rom_memory[21629] = 3'b110;
        rom_memory[21630] = 3'b111;
        rom_memory[21631] = 3'b111;
        rom_memory[21632] = 3'b111;
        rom_memory[21633] = 3'b111;
        rom_memory[21634] = 3'b111;
        rom_memory[21635] = 3'b111;
        rom_memory[21636] = 3'b111;
        rom_memory[21637] = 3'b111;
        rom_memory[21638] = 3'b111;
        rom_memory[21639] = 3'b111;
        rom_memory[21640] = 3'b111;
        rom_memory[21641] = 3'b111;
        rom_memory[21642] = 3'b111;
        rom_memory[21643] = 3'b111;
        rom_memory[21644] = 3'b111;
        rom_memory[21645] = 3'b111;
        rom_memory[21646] = 3'b111;
        rom_memory[21647] = 3'b110;
        rom_memory[21648] = 3'b110;
        rom_memory[21649] = 3'b100;
        rom_memory[21650] = 3'b110;
        rom_memory[21651] = 3'b110;
        rom_memory[21652] = 3'b110;
        rom_memory[21653] = 3'b110;
        rom_memory[21654] = 3'b110;
        rom_memory[21655] = 3'b110;
        rom_memory[21656] = 3'b100;
        rom_memory[21657] = 3'b100;
        rom_memory[21658] = 3'b100;
        rom_memory[21659] = 3'b100;
        rom_memory[21660] = 3'b100;
        rom_memory[21661] = 3'b110;
        rom_memory[21662] = 3'b100;
        rom_memory[21663] = 3'b100;
        rom_memory[21664] = 3'b110;
        rom_memory[21665] = 3'b110;
        rom_memory[21666] = 3'b110;
        rom_memory[21667] = 3'b110;
        rom_memory[21668] = 3'b110;
        rom_memory[21669] = 3'b110;
        rom_memory[21670] = 3'b110;
        rom_memory[21671] = 3'b110;
        rom_memory[21672] = 3'b110;
        rom_memory[21673] = 3'b110;
        rom_memory[21674] = 3'b110;
        rom_memory[21675] = 3'b110;
        rom_memory[21676] = 3'b110;
        rom_memory[21677] = 3'b110;
        rom_memory[21678] = 3'b110;
        rom_memory[21679] = 3'b110;
        rom_memory[21680] = 3'b110;
        rom_memory[21681] = 3'b110;
        rom_memory[21682] = 3'b110;
        rom_memory[21683] = 3'b110;
        rom_memory[21684] = 3'b110;
        rom_memory[21685] = 3'b110;
        rom_memory[21686] = 3'b110;
        rom_memory[21687] = 3'b110;
        rom_memory[21688] = 3'b110;
        rom_memory[21689] = 3'b110;
        rom_memory[21690] = 3'b110;
        rom_memory[21691] = 3'b110;
        rom_memory[21692] = 3'b110;
        rom_memory[21693] = 3'b110;
        rom_memory[21694] = 3'b110;
        rom_memory[21695] = 3'b110;
        rom_memory[21696] = 3'b110;
        rom_memory[21697] = 3'b110;
        rom_memory[21698] = 3'b111;
        rom_memory[21699] = 3'b111;
        rom_memory[21700] = 3'b111;
        rom_memory[21701] = 3'b111;
        rom_memory[21702] = 3'b111;
        rom_memory[21703] = 3'b111;
        rom_memory[21704] = 3'b111;
        rom_memory[21705] = 3'b100;
        rom_memory[21706] = 3'b000;
        rom_memory[21707] = 3'b000;
        rom_memory[21708] = 3'b000;
        rom_memory[21709] = 3'b000;
        rom_memory[21710] = 3'b000;
        rom_memory[21711] = 3'b000;
        rom_memory[21712] = 3'b000;
        rom_memory[21713] = 3'b000;
        rom_memory[21714] = 3'b100;
        rom_memory[21715] = 3'b000;
        rom_memory[21716] = 3'b110;
        rom_memory[21717] = 3'b100;
        rom_memory[21718] = 3'b110;
        rom_memory[21719] = 3'b110;
        rom_memory[21720] = 3'b110;
        rom_memory[21721] = 3'b110;
        rom_memory[21722] = 3'b110;
        rom_memory[21723] = 3'b110;
        rom_memory[21724] = 3'b110;
        rom_memory[21725] = 3'b111;
        rom_memory[21726] = 3'b111;
        rom_memory[21727] = 3'b110;
        rom_memory[21728] = 3'b110;
        rom_memory[21729] = 3'b110;
        rom_memory[21730] = 3'b110;
        rom_memory[21731] = 3'b110;
        rom_memory[21732] = 3'b110;
        rom_memory[21733] = 3'b110;
        rom_memory[21734] = 3'b110;
        rom_memory[21735] = 3'b110;
        rom_memory[21736] = 3'b110;
        rom_memory[21737] = 3'b110;
        rom_memory[21738] = 3'b110;
        rom_memory[21739] = 3'b110;
        rom_memory[21740] = 3'b110;
        rom_memory[21741] = 3'b110;
        rom_memory[21742] = 3'b110;
        rom_memory[21743] = 3'b110;
        rom_memory[21744] = 3'b110;
        rom_memory[21745] = 3'b110;
        rom_memory[21746] = 3'b110;
        rom_memory[21747] = 3'b110;
        rom_memory[21748] = 3'b111;
        rom_memory[21749] = 3'b110;
        rom_memory[21750] = 3'b111;
        rom_memory[21751] = 3'b111;
        rom_memory[21752] = 3'b111;
        rom_memory[21753] = 3'b111;
        rom_memory[21754] = 3'b111;
        rom_memory[21755] = 3'b111;
        rom_memory[21756] = 3'b111;
        rom_memory[21757] = 3'b111;
        rom_memory[21758] = 3'b111;
        rom_memory[21759] = 3'b111;
        rom_memory[21760] = 3'b111;
        rom_memory[21761] = 3'b111;
        rom_memory[21762] = 3'b111;
        rom_memory[21763] = 3'b111;
        rom_memory[21764] = 3'b111;
        rom_memory[21765] = 3'b111;
        rom_memory[21766] = 3'b111;
        rom_memory[21767] = 3'b111;
        rom_memory[21768] = 3'b111;
        rom_memory[21769] = 3'b111;
        rom_memory[21770] = 3'b111;
        rom_memory[21771] = 3'b111;
        rom_memory[21772] = 3'b111;
        rom_memory[21773] = 3'b111;
        rom_memory[21774] = 3'b111;
        rom_memory[21775] = 3'b111;
        rom_memory[21776] = 3'b111;
        rom_memory[21777] = 3'b111;
        rom_memory[21778] = 3'b111;
        rom_memory[21779] = 3'b111;
        rom_memory[21780] = 3'b111;
        rom_memory[21781] = 3'b111;
        rom_memory[21782] = 3'b111;
        rom_memory[21783] = 3'b111;
        rom_memory[21784] = 3'b111;
        rom_memory[21785] = 3'b111;
        rom_memory[21786] = 3'b111;
        rom_memory[21787] = 3'b111;
        rom_memory[21788] = 3'b111;
        rom_memory[21789] = 3'b111;
        rom_memory[21790] = 3'b111;
        rom_memory[21791] = 3'b111;
        rom_memory[21792] = 3'b110;
        rom_memory[21793] = 3'b110;
        rom_memory[21794] = 3'b110;
        rom_memory[21795] = 3'b110;
        rom_memory[21796] = 3'b110;
        rom_memory[21797] = 3'b110;
        rom_memory[21798] = 3'b110;
        rom_memory[21799] = 3'b110;
        rom_memory[21800] = 3'b110;
        rom_memory[21801] = 3'b111;
        rom_memory[21802] = 3'b110;
        rom_memory[21803] = 3'b110;
        rom_memory[21804] = 3'b111;
        rom_memory[21805] = 3'b110;
        rom_memory[21806] = 3'b110;
        rom_memory[21807] = 3'b110;
        rom_memory[21808] = 3'b110;
        rom_memory[21809] = 3'b110;
        rom_memory[21810] = 3'b110;
        rom_memory[21811] = 3'b110;
        rom_memory[21812] = 3'b110;
        rom_memory[21813] = 3'b110;
        rom_memory[21814] = 3'b110;
        rom_memory[21815] = 3'b110;
        rom_memory[21816] = 3'b110;
        rom_memory[21817] = 3'b110;
        rom_memory[21818] = 3'b110;
        rom_memory[21819] = 3'b110;
        rom_memory[21820] = 3'b110;
        rom_memory[21821] = 3'b110;
        rom_memory[21822] = 3'b110;
        rom_memory[21823] = 3'b110;
        rom_memory[21824] = 3'b110;
        rom_memory[21825] = 3'b110;
        rom_memory[21826] = 3'b110;
        rom_memory[21827] = 3'b110;
        rom_memory[21828] = 3'b110;
        rom_memory[21829] = 3'b110;
        rom_memory[21830] = 3'b110;
        rom_memory[21831] = 3'b110;
        rom_memory[21832] = 3'b110;
        rom_memory[21833] = 3'b110;
        rom_memory[21834] = 3'b110;
        rom_memory[21835] = 3'b110;
        rom_memory[21836] = 3'b110;
        rom_memory[21837] = 3'b110;
        rom_memory[21838] = 3'b110;
        rom_memory[21839] = 3'b110;
        rom_memory[21840] = 3'b110;
        rom_memory[21841] = 3'b110;
        rom_memory[21842] = 3'b110;
        rom_memory[21843] = 3'b110;
        rom_memory[21844] = 3'b110;
        rom_memory[21845] = 3'b110;
        rom_memory[21846] = 3'b110;
        rom_memory[21847] = 3'b110;
        rom_memory[21848] = 3'b110;
        rom_memory[21849] = 3'b110;
        rom_memory[21850] = 3'b110;
        rom_memory[21851] = 3'b110;
        rom_memory[21852] = 3'b110;
        rom_memory[21853] = 3'b110;
        rom_memory[21854] = 3'b110;
        rom_memory[21855] = 3'b110;
        rom_memory[21856] = 3'b110;
        rom_memory[21857] = 3'b110;
        rom_memory[21858] = 3'b110;
        rom_memory[21859] = 3'b110;
        rom_memory[21860] = 3'b110;
        rom_memory[21861] = 3'b110;
        rom_memory[21862] = 3'b110;
        rom_memory[21863] = 3'b110;
        rom_memory[21864] = 3'b110;
        rom_memory[21865] = 3'b110;
        rom_memory[21866] = 3'b110;
        rom_memory[21867] = 3'b110;
        rom_memory[21868] = 3'b110;
        rom_memory[21869] = 3'b110;
        rom_memory[21870] = 3'b111;
        rom_memory[21871] = 3'b111;
        rom_memory[21872] = 3'b111;
        rom_memory[21873] = 3'b111;
        rom_memory[21874] = 3'b111;
        rom_memory[21875] = 3'b111;
        rom_memory[21876] = 3'b111;
        rom_memory[21877] = 3'b111;
        rom_memory[21878] = 3'b111;
        rom_memory[21879] = 3'b111;
        rom_memory[21880] = 3'b111;
        rom_memory[21881] = 3'b111;
        rom_memory[21882] = 3'b111;
        rom_memory[21883] = 3'b111;
        rom_memory[21884] = 3'b111;
        rom_memory[21885] = 3'b111;
        rom_memory[21886] = 3'b111;
        rom_memory[21887] = 3'b111;
        rom_memory[21888] = 3'b110;
        rom_memory[21889] = 3'b100;
        rom_memory[21890] = 3'b110;
        rom_memory[21891] = 3'b110;
        rom_memory[21892] = 3'b110;
        rom_memory[21893] = 3'b110;
        rom_memory[21894] = 3'b110;
        rom_memory[21895] = 3'b110;
        rom_memory[21896] = 3'b110;
        rom_memory[21897] = 3'b100;
        rom_memory[21898] = 3'b100;
        rom_memory[21899] = 3'b100;
        rom_memory[21900] = 3'b100;
        rom_memory[21901] = 3'b110;
        rom_memory[21902] = 3'b100;
        rom_memory[21903] = 3'b100;
        rom_memory[21904] = 3'b100;
        rom_memory[21905] = 3'b110;
        rom_memory[21906] = 3'b110;
        rom_memory[21907] = 3'b110;
        rom_memory[21908] = 3'b110;
        rom_memory[21909] = 3'b110;
        rom_memory[21910] = 3'b110;
        rom_memory[21911] = 3'b110;
        rom_memory[21912] = 3'b110;
        rom_memory[21913] = 3'b110;
        rom_memory[21914] = 3'b110;
        rom_memory[21915] = 3'b110;
        rom_memory[21916] = 3'b110;
        rom_memory[21917] = 3'b110;
        rom_memory[21918] = 3'b110;
        rom_memory[21919] = 3'b110;
        rom_memory[21920] = 3'b110;
        rom_memory[21921] = 3'b110;
        rom_memory[21922] = 3'b110;
        rom_memory[21923] = 3'b110;
        rom_memory[21924] = 3'b110;
        rom_memory[21925] = 3'b110;
        rom_memory[21926] = 3'b110;
        rom_memory[21927] = 3'b110;
        rom_memory[21928] = 3'b110;
        rom_memory[21929] = 3'b110;
        rom_memory[21930] = 3'b110;
        rom_memory[21931] = 3'b110;
        rom_memory[21932] = 3'b110;
        rom_memory[21933] = 3'b110;
        rom_memory[21934] = 3'b110;
        rom_memory[21935] = 3'b110;
        rom_memory[21936] = 3'b110;
        rom_memory[21937] = 3'b110;
        rom_memory[21938] = 3'b110;
        rom_memory[21939] = 3'b111;
        rom_memory[21940] = 3'b111;
        rom_memory[21941] = 3'b111;
        rom_memory[21942] = 3'b111;
        rom_memory[21943] = 3'b111;
        rom_memory[21944] = 3'b111;
        rom_memory[21945] = 3'b111;
        rom_memory[21946] = 3'b110;
        rom_memory[21947] = 3'b000;
        rom_memory[21948] = 3'b000;
        rom_memory[21949] = 3'b000;
        rom_memory[21950] = 3'b000;
        rom_memory[21951] = 3'b000;
        rom_memory[21952] = 3'b000;
        rom_memory[21953] = 3'b000;
        rom_memory[21954] = 3'b000;
        rom_memory[21955] = 3'b100;
        rom_memory[21956] = 3'b000;
        rom_memory[21957] = 3'b110;
        rom_memory[21958] = 3'b100;
        rom_memory[21959] = 3'b110;
        rom_memory[21960] = 3'b110;
        rom_memory[21961] = 3'b110;
        rom_memory[21962] = 3'b110;
        rom_memory[21963] = 3'b110;
        rom_memory[21964] = 3'b110;
        rom_memory[21965] = 3'b111;
        rom_memory[21966] = 3'b111;
        rom_memory[21967] = 3'b111;
        rom_memory[21968] = 3'b110;
        rom_memory[21969] = 3'b110;
        rom_memory[21970] = 3'b110;
        rom_memory[21971] = 3'b110;
        rom_memory[21972] = 3'b110;
        rom_memory[21973] = 3'b110;
        rom_memory[21974] = 3'b110;
        rom_memory[21975] = 3'b110;
        rom_memory[21976] = 3'b110;
        rom_memory[21977] = 3'b110;
        rom_memory[21978] = 3'b110;
        rom_memory[21979] = 3'b110;
        rom_memory[21980] = 3'b110;
        rom_memory[21981] = 3'b110;
        rom_memory[21982] = 3'b110;
        rom_memory[21983] = 3'b110;
        rom_memory[21984] = 3'b110;
        rom_memory[21985] = 3'b110;
        rom_memory[21986] = 3'b110;
        rom_memory[21987] = 3'b110;
        rom_memory[21988] = 3'b111;
        rom_memory[21989] = 3'b111;
        rom_memory[21990] = 3'b111;
        rom_memory[21991] = 3'b110;
        rom_memory[21992] = 3'b111;
        rom_memory[21993] = 3'b111;
        rom_memory[21994] = 3'b111;
        rom_memory[21995] = 3'b111;
        rom_memory[21996] = 3'b111;
        rom_memory[21997] = 3'b111;
        rom_memory[21998] = 3'b111;
        rom_memory[21999] = 3'b111;
        rom_memory[22000] = 3'b111;
        rom_memory[22001] = 3'b111;
        rom_memory[22002] = 3'b111;
        rom_memory[22003] = 3'b111;
        rom_memory[22004] = 3'b111;
        rom_memory[22005] = 3'b111;
        rom_memory[22006] = 3'b111;
        rom_memory[22007] = 3'b111;
        rom_memory[22008] = 3'b111;
        rom_memory[22009] = 3'b111;
        rom_memory[22010] = 3'b111;
        rom_memory[22011] = 3'b111;
        rom_memory[22012] = 3'b111;
        rom_memory[22013] = 3'b111;
        rom_memory[22014] = 3'b111;
        rom_memory[22015] = 3'b111;
        rom_memory[22016] = 3'b111;
        rom_memory[22017] = 3'b111;
        rom_memory[22018] = 3'b111;
        rom_memory[22019] = 3'b111;
        rom_memory[22020] = 3'b111;
        rom_memory[22021] = 3'b111;
        rom_memory[22022] = 3'b111;
        rom_memory[22023] = 3'b111;
        rom_memory[22024] = 3'b111;
        rom_memory[22025] = 3'b111;
        rom_memory[22026] = 3'b111;
        rom_memory[22027] = 3'b111;
        rom_memory[22028] = 3'b111;
        rom_memory[22029] = 3'b111;
        rom_memory[22030] = 3'b111;
        rom_memory[22031] = 3'b111;
        rom_memory[22032] = 3'b111;
        rom_memory[22033] = 3'b111;
        rom_memory[22034] = 3'b111;
        rom_memory[22035] = 3'b110;
        rom_memory[22036] = 3'b111;
        rom_memory[22037] = 3'b111;
        rom_memory[22038] = 3'b110;
        rom_memory[22039] = 3'b110;
        rom_memory[22040] = 3'b110;
        rom_memory[22041] = 3'b110;
        rom_memory[22042] = 3'b110;
        rom_memory[22043] = 3'b110;
        rom_memory[22044] = 3'b111;
        rom_memory[22045] = 3'b111;
        rom_memory[22046] = 3'b110;
        rom_memory[22047] = 3'b110;
        rom_memory[22048] = 3'b110;
        rom_memory[22049] = 3'b110;
        rom_memory[22050] = 3'b111;
        rom_memory[22051] = 3'b110;
        rom_memory[22052] = 3'b110;
        rom_memory[22053] = 3'b110;
        rom_memory[22054] = 3'b110;
        rom_memory[22055] = 3'b110;
        rom_memory[22056] = 3'b111;
        rom_memory[22057] = 3'b110;
        rom_memory[22058] = 3'b110;
        rom_memory[22059] = 3'b111;
        rom_memory[22060] = 3'b110;
        rom_memory[22061] = 3'b110;
        rom_memory[22062] = 3'b110;
        rom_memory[22063] = 3'b110;
        rom_memory[22064] = 3'b110;
        rom_memory[22065] = 3'b110;
        rom_memory[22066] = 3'b110;
        rom_memory[22067] = 3'b110;
        rom_memory[22068] = 3'b110;
        rom_memory[22069] = 3'b110;
        rom_memory[22070] = 3'b110;
        rom_memory[22071] = 3'b110;
        rom_memory[22072] = 3'b110;
        rom_memory[22073] = 3'b110;
        rom_memory[22074] = 3'b110;
        rom_memory[22075] = 3'b110;
        rom_memory[22076] = 3'b110;
        rom_memory[22077] = 3'b110;
        rom_memory[22078] = 3'b110;
        rom_memory[22079] = 3'b110;
        rom_memory[22080] = 3'b110;
        rom_memory[22081] = 3'b110;
        rom_memory[22082] = 3'b110;
        rom_memory[22083] = 3'b110;
        rom_memory[22084] = 3'b110;
        rom_memory[22085] = 3'b110;
        rom_memory[22086] = 3'b110;
        rom_memory[22087] = 3'b110;
        rom_memory[22088] = 3'b110;
        rom_memory[22089] = 3'b110;
        rom_memory[22090] = 3'b110;
        rom_memory[22091] = 3'b110;
        rom_memory[22092] = 3'b110;
        rom_memory[22093] = 3'b110;
        rom_memory[22094] = 3'b110;
        rom_memory[22095] = 3'b110;
        rom_memory[22096] = 3'b110;
        rom_memory[22097] = 3'b110;
        rom_memory[22098] = 3'b110;
        rom_memory[22099] = 3'b110;
        rom_memory[22100] = 3'b110;
        rom_memory[22101] = 3'b110;
        rom_memory[22102] = 3'b110;
        rom_memory[22103] = 3'b110;
        rom_memory[22104] = 3'b110;
        rom_memory[22105] = 3'b110;
        rom_memory[22106] = 3'b110;
        rom_memory[22107] = 3'b110;
        rom_memory[22108] = 3'b110;
        rom_memory[22109] = 3'b111;
        rom_memory[22110] = 3'b111;
        rom_memory[22111] = 3'b111;
        rom_memory[22112] = 3'b111;
        rom_memory[22113] = 3'b111;
        rom_memory[22114] = 3'b111;
        rom_memory[22115] = 3'b111;
        rom_memory[22116] = 3'b111;
        rom_memory[22117] = 3'b111;
        rom_memory[22118] = 3'b111;
        rom_memory[22119] = 3'b111;
        rom_memory[22120] = 3'b111;
        rom_memory[22121] = 3'b111;
        rom_memory[22122] = 3'b111;
        rom_memory[22123] = 3'b111;
        rom_memory[22124] = 3'b111;
        rom_memory[22125] = 3'b111;
        rom_memory[22126] = 3'b111;
        rom_memory[22127] = 3'b111;
        rom_memory[22128] = 3'b110;
        rom_memory[22129] = 3'b100;
        rom_memory[22130] = 3'b100;
        rom_memory[22131] = 3'b100;
        rom_memory[22132] = 3'b110;
        rom_memory[22133] = 3'b110;
        rom_memory[22134] = 3'b110;
        rom_memory[22135] = 3'b110;
        rom_memory[22136] = 3'b110;
        rom_memory[22137] = 3'b100;
        rom_memory[22138] = 3'b100;
        rom_memory[22139] = 3'b100;
        rom_memory[22140] = 3'b100;
        rom_memory[22141] = 3'b110;
        rom_memory[22142] = 3'b110;
        rom_memory[22143] = 3'b100;
        rom_memory[22144] = 3'b100;
        rom_memory[22145] = 3'b110;
        rom_memory[22146] = 3'b110;
        rom_memory[22147] = 3'b110;
        rom_memory[22148] = 3'b110;
        rom_memory[22149] = 3'b110;
        rom_memory[22150] = 3'b110;
        rom_memory[22151] = 3'b110;
        rom_memory[22152] = 3'b110;
        rom_memory[22153] = 3'b110;
        rom_memory[22154] = 3'b110;
        rom_memory[22155] = 3'b110;
        rom_memory[22156] = 3'b110;
        rom_memory[22157] = 3'b110;
        rom_memory[22158] = 3'b110;
        rom_memory[22159] = 3'b110;
        rom_memory[22160] = 3'b110;
        rom_memory[22161] = 3'b110;
        rom_memory[22162] = 3'b110;
        rom_memory[22163] = 3'b110;
        rom_memory[22164] = 3'b110;
        rom_memory[22165] = 3'b110;
        rom_memory[22166] = 3'b110;
        rom_memory[22167] = 3'b110;
        rom_memory[22168] = 3'b110;
        rom_memory[22169] = 3'b110;
        rom_memory[22170] = 3'b110;
        rom_memory[22171] = 3'b110;
        rom_memory[22172] = 3'b110;
        rom_memory[22173] = 3'b110;
        rom_memory[22174] = 3'b110;
        rom_memory[22175] = 3'b110;
        rom_memory[22176] = 3'b110;
        rom_memory[22177] = 3'b110;
        rom_memory[22178] = 3'b110;
        rom_memory[22179] = 3'b110;
        rom_memory[22180] = 3'b111;
        rom_memory[22181] = 3'b111;
        rom_memory[22182] = 3'b111;
        rom_memory[22183] = 3'b111;
        rom_memory[22184] = 3'b111;
        rom_memory[22185] = 3'b111;
        rom_memory[22186] = 3'b111;
        rom_memory[22187] = 3'b110;
        rom_memory[22188] = 3'b000;
        rom_memory[22189] = 3'b000;
        rom_memory[22190] = 3'b000;
        rom_memory[22191] = 3'b000;
        rom_memory[22192] = 3'b000;
        rom_memory[22193] = 3'b000;
        rom_memory[22194] = 3'b000;
        rom_memory[22195] = 3'b000;
        rom_memory[22196] = 3'b100;
        rom_memory[22197] = 3'b100;
        rom_memory[22198] = 3'b110;
        rom_memory[22199] = 3'b000;
        rom_memory[22200] = 3'b100;
        rom_memory[22201] = 3'b110;
        rom_memory[22202] = 3'b110;
        rom_memory[22203] = 3'b110;
        rom_memory[22204] = 3'b110;
        rom_memory[22205] = 3'b111;
        rom_memory[22206] = 3'b110;
        rom_memory[22207] = 3'b111;
        rom_memory[22208] = 3'b110;
        rom_memory[22209] = 3'b110;
        rom_memory[22210] = 3'b110;
        rom_memory[22211] = 3'b110;
        rom_memory[22212] = 3'b110;
        rom_memory[22213] = 3'b110;
        rom_memory[22214] = 3'b110;
        rom_memory[22215] = 3'b110;
        rom_memory[22216] = 3'b110;
        rom_memory[22217] = 3'b110;
        rom_memory[22218] = 3'b110;
        rom_memory[22219] = 3'b110;
        rom_memory[22220] = 3'b110;
        rom_memory[22221] = 3'b110;
        rom_memory[22222] = 3'b110;
        rom_memory[22223] = 3'b110;
        rom_memory[22224] = 3'b110;
        rom_memory[22225] = 3'b110;
        rom_memory[22226] = 3'b110;
        rom_memory[22227] = 3'b110;
        rom_memory[22228] = 3'b110;
        rom_memory[22229] = 3'b110;
        rom_memory[22230] = 3'b110;
        rom_memory[22231] = 3'b110;
        rom_memory[22232] = 3'b111;
        rom_memory[22233] = 3'b111;
        rom_memory[22234] = 3'b110;
        rom_memory[22235] = 3'b111;
        rom_memory[22236] = 3'b111;
        rom_memory[22237] = 3'b111;
        rom_memory[22238] = 3'b111;
        rom_memory[22239] = 3'b111;
        rom_memory[22240] = 3'b111;
        rom_memory[22241] = 3'b111;
        rom_memory[22242] = 3'b111;
        rom_memory[22243] = 3'b111;
        rom_memory[22244] = 3'b111;
        rom_memory[22245] = 3'b111;
        rom_memory[22246] = 3'b111;
        rom_memory[22247] = 3'b111;
        rom_memory[22248] = 3'b111;
        rom_memory[22249] = 3'b111;
        rom_memory[22250] = 3'b111;
        rom_memory[22251] = 3'b111;
        rom_memory[22252] = 3'b111;
        rom_memory[22253] = 3'b111;
        rom_memory[22254] = 3'b111;
        rom_memory[22255] = 3'b111;
        rom_memory[22256] = 3'b111;
        rom_memory[22257] = 3'b111;
        rom_memory[22258] = 3'b111;
        rom_memory[22259] = 3'b111;
        rom_memory[22260] = 3'b111;
        rom_memory[22261] = 3'b111;
        rom_memory[22262] = 3'b111;
        rom_memory[22263] = 3'b111;
        rom_memory[22264] = 3'b111;
        rom_memory[22265] = 3'b111;
        rom_memory[22266] = 3'b111;
        rom_memory[22267] = 3'b111;
        rom_memory[22268] = 3'b110;
        rom_memory[22269] = 3'b111;
        rom_memory[22270] = 3'b110;
        rom_memory[22271] = 3'b111;
        rom_memory[22272] = 3'b111;
        rom_memory[22273] = 3'b110;
        rom_memory[22274] = 3'b110;
        rom_memory[22275] = 3'b110;
        rom_memory[22276] = 3'b110;
        rom_memory[22277] = 3'b110;
        rom_memory[22278] = 3'b110;
        rom_memory[22279] = 3'b110;
        rom_memory[22280] = 3'b110;
        rom_memory[22281] = 3'b110;
        rom_memory[22282] = 3'b111;
        rom_memory[22283] = 3'b111;
        rom_memory[22284] = 3'b111;
        rom_memory[22285] = 3'b111;
        rom_memory[22286] = 3'b111;
        rom_memory[22287] = 3'b111;
        rom_memory[22288] = 3'b111;
        rom_memory[22289] = 3'b110;
        rom_memory[22290] = 3'b111;
        rom_memory[22291] = 3'b110;
        rom_memory[22292] = 3'b110;
        rom_memory[22293] = 3'b111;
        rom_memory[22294] = 3'b111;
        rom_memory[22295] = 3'b110;
        rom_memory[22296] = 3'b110;
        rom_memory[22297] = 3'b110;
        rom_memory[22298] = 3'b110;
        rom_memory[22299] = 3'b111;
        rom_memory[22300] = 3'b111;
        rom_memory[22301] = 3'b111;
        rom_memory[22302] = 3'b111;
        rom_memory[22303] = 3'b110;
        rom_memory[22304] = 3'b111;
        rom_memory[22305] = 3'b110;
        rom_memory[22306] = 3'b110;
        rom_memory[22307] = 3'b110;
        rom_memory[22308] = 3'b111;
        rom_memory[22309] = 3'b111;
        rom_memory[22310] = 3'b110;
        rom_memory[22311] = 3'b111;
        rom_memory[22312] = 3'b110;
        rom_memory[22313] = 3'b110;
        rom_memory[22314] = 3'b110;
        rom_memory[22315] = 3'b110;
        rom_memory[22316] = 3'b110;
        rom_memory[22317] = 3'b110;
        rom_memory[22318] = 3'b110;
        rom_memory[22319] = 3'b110;
        rom_memory[22320] = 3'b110;
        rom_memory[22321] = 3'b110;
        rom_memory[22322] = 3'b110;
        rom_memory[22323] = 3'b110;
        rom_memory[22324] = 3'b110;
        rom_memory[22325] = 3'b110;
        rom_memory[22326] = 3'b110;
        rom_memory[22327] = 3'b110;
        rom_memory[22328] = 3'b110;
        rom_memory[22329] = 3'b110;
        rom_memory[22330] = 3'b110;
        rom_memory[22331] = 3'b110;
        rom_memory[22332] = 3'b110;
        rom_memory[22333] = 3'b110;
        rom_memory[22334] = 3'b110;
        rom_memory[22335] = 3'b110;
        rom_memory[22336] = 3'b110;
        rom_memory[22337] = 3'b110;
        rom_memory[22338] = 3'b110;
        rom_memory[22339] = 3'b110;
        rom_memory[22340] = 3'b110;
        rom_memory[22341] = 3'b110;
        rom_memory[22342] = 3'b110;
        rom_memory[22343] = 3'b110;
        rom_memory[22344] = 3'b110;
        rom_memory[22345] = 3'b110;
        rom_memory[22346] = 3'b110;
        rom_memory[22347] = 3'b110;
        rom_memory[22348] = 3'b110;
        rom_memory[22349] = 3'b111;
        rom_memory[22350] = 3'b111;
        rom_memory[22351] = 3'b111;
        rom_memory[22352] = 3'b111;
        rom_memory[22353] = 3'b111;
        rom_memory[22354] = 3'b111;
        rom_memory[22355] = 3'b111;
        rom_memory[22356] = 3'b111;
        rom_memory[22357] = 3'b111;
        rom_memory[22358] = 3'b111;
        rom_memory[22359] = 3'b111;
        rom_memory[22360] = 3'b111;
        rom_memory[22361] = 3'b111;
        rom_memory[22362] = 3'b111;
        rom_memory[22363] = 3'b111;
        rom_memory[22364] = 3'b111;
        rom_memory[22365] = 3'b111;
        rom_memory[22366] = 3'b111;
        rom_memory[22367] = 3'b111;
        rom_memory[22368] = 3'b110;
        rom_memory[22369] = 3'b100;
        rom_memory[22370] = 3'b100;
        rom_memory[22371] = 3'b100;
        rom_memory[22372] = 3'b100;
        rom_memory[22373] = 3'b110;
        rom_memory[22374] = 3'b110;
        rom_memory[22375] = 3'b110;
        rom_memory[22376] = 3'b110;
        rom_memory[22377] = 3'b100;
        rom_memory[22378] = 3'b100;
        rom_memory[22379] = 3'b100;
        rom_memory[22380] = 3'b100;
        rom_memory[22381] = 3'b110;
        rom_memory[22382] = 3'b110;
        rom_memory[22383] = 3'b110;
        rom_memory[22384] = 3'b110;
        rom_memory[22385] = 3'b110;
        rom_memory[22386] = 3'b110;
        rom_memory[22387] = 3'b110;
        rom_memory[22388] = 3'b110;
        rom_memory[22389] = 3'b110;
        rom_memory[22390] = 3'b110;
        rom_memory[22391] = 3'b110;
        rom_memory[22392] = 3'b110;
        rom_memory[22393] = 3'b110;
        rom_memory[22394] = 3'b110;
        rom_memory[22395] = 3'b110;
        rom_memory[22396] = 3'b110;
        rom_memory[22397] = 3'b110;
        rom_memory[22398] = 3'b110;
        rom_memory[22399] = 3'b110;
        rom_memory[22400] = 3'b110;
        rom_memory[22401] = 3'b110;
        rom_memory[22402] = 3'b110;
        rom_memory[22403] = 3'b110;
        rom_memory[22404] = 3'b110;
        rom_memory[22405] = 3'b110;
        rom_memory[22406] = 3'b110;
        rom_memory[22407] = 3'b110;
        rom_memory[22408] = 3'b110;
        rom_memory[22409] = 3'b110;
        rom_memory[22410] = 3'b110;
        rom_memory[22411] = 3'b110;
        rom_memory[22412] = 3'b110;
        rom_memory[22413] = 3'b110;
        rom_memory[22414] = 3'b110;
        rom_memory[22415] = 3'b110;
        rom_memory[22416] = 3'b110;
        rom_memory[22417] = 3'b110;
        rom_memory[22418] = 3'b110;
        rom_memory[22419] = 3'b110;
        rom_memory[22420] = 3'b111;
        rom_memory[22421] = 3'b111;
        rom_memory[22422] = 3'b111;
        rom_memory[22423] = 3'b111;
        rom_memory[22424] = 3'b111;
        rom_memory[22425] = 3'b111;
        rom_memory[22426] = 3'b111;
        rom_memory[22427] = 3'b111;
        rom_memory[22428] = 3'b111;
        rom_memory[22429] = 3'b000;
        rom_memory[22430] = 3'b000;
        rom_memory[22431] = 3'b000;
        rom_memory[22432] = 3'b000;
        rom_memory[22433] = 3'b000;
        rom_memory[22434] = 3'b000;
        rom_memory[22435] = 3'b000;
        rom_memory[22436] = 3'b000;
        rom_memory[22437] = 3'b100;
        rom_memory[22438] = 3'b000;
        rom_memory[22439] = 3'b110;
        rom_memory[22440] = 3'b000;
        rom_memory[22441] = 3'b100;
        rom_memory[22442] = 3'b110;
        rom_memory[22443] = 3'b110;
        rom_memory[22444] = 3'b110;
        rom_memory[22445] = 3'b111;
        rom_memory[22446] = 3'b111;
        rom_memory[22447] = 3'b111;
        rom_memory[22448] = 3'b111;
        rom_memory[22449] = 3'b110;
        rom_memory[22450] = 3'b110;
        rom_memory[22451] = 3'b110;
        rom_memory[22452] = 3'b110;
        rom_memory[22453] = 3'b110;
        rom_memory[22454] = 3'b110;
        rom_memory[22455] = 3'b110;
        rom_memory[22456] = 3'b110;
        rom_memory[22457] = 3'b110;
        rom_memory[22458] = 3'b110;
        rom_memory[22459] = 3'b110;
        rom_memory[22460] = 3'b110;
        rom_memory[22461] = 3'b110;
        rom_memory[22462] = 3'b110;
        rom_memory[22463] = 3'b110;
        rom_memory[22464] = 3'b110;
        rom_memory[22465] = 3'b110;
        rom_memory[22466] = 3'b110;
        rom_memory[22467] = 3'b110;
        rom_memory[22468] = 3'b110;
        rom_memory[22469] = 3'b110;
        rom_memory[22470] = 3'b110;
        rom_memory[22471] = 3'b110;
        rom_memory[22472] = 3'b111;
        rom_memory[22473] = 3'b111;
        rom_memory[22474] = 3'b111;
        rom_memory[22475] = 3'b111;
        rom_memory[22476] = 3'b111;
        rom_memory[22477] = 3'b111;
        rom_memory[22478] = 3'b111;
        rom_memory[22479] = 3'b111;
        rom_memory[22480] = 3'b111;
        rom_memory[22481] = 3'b111;
        rom_memory[22482] = 3'b111;
        rom_memory[22483] = 3'b111;
        rom_memory[22484] = 3'b111;
        rom_memory[22485] = 3'b111;
        rom_memory[22486] = 3'b111;
        rom_memory[22487] = 3'b111;
        rom_memory[22488] = 3'b111;
        rom_memory[22489] = 3'b111;
        rom_memory[22490] = 3'b111;
        rom_memory[22491] = 3'b111;
        rom_memory[22492] = 3'b111;
        rom_memory[22493] = 3'b111;
        rom_memory[22494] = 3'b111;
        rom_memory[22495] = 3'b111;
        rom_memory[22496] = 3'b111;
        rom_memory[22497] = 3'b111;
        rom_memory[22498] = 3'b111;
        rom_memory[22499] = 3'b111;
        rom_memory[22500] = 3'b111;
        rom_memory[22501] = 3'b111;
        rom_memory[22502] = 3'b111;
        rom_memory[22503] = 3'b111;
        rom_memory[22504] = 3'b111;
        rom_memory[22505] = 3'b111;
        rom_memory[22506] = 3'b111;
        rom_memory[22507] = 3'b111;
        rom_memory[22508] = 3'b110;
        rom_memory[22509] = 3'b111;
        rom_memory[22510] = 3'b111;
        rom_memory[22511] = 3'b111;
        rom_memory[22512] = 3'b110;
        rom_memory[22513] = 3'b110;
        rom_memory[22514] = 3'b110;
        rom_memory[22515] = 3'b110;
        rom_memory[22516] = 3'b110;
        rom_memory[22517] = 3'b110;
        rom_memory[22518] = 3'b111;
        rom_memory[22519] = 3'b111;
        rom_memory[22520] = 3'b111;
        rom_memory[22521] = 3'b111;
        rom_memory[22522] = 3'b111;
        rom_memory[22523] = 3'b111;
        rom_memory[22524] = 3'b111;
        rom_memory[22525] = 3'b111;
        rom_memory[22526] = 3'b111;
        rom_memory[22527] = 3'b111;
        rom_memory[22528] = 3'b111;
        rom_memory[22529] = 3'b111;
        rom_memory[22530] = 3'b111;
        rom_memory[22531] = 3'b110;
        rom_memory[22532] = 3'b111;
        rom_memory[22533] = 3'b111;
        rom_memory[22534] = 3'b110;
        rom_memory[22535] = 3'b110;
        rom_memory[22536] = 3'b110;
        rom_memory[22537] = 3'b110;
        rom_memory[22538] = 3'b111;
        rom_memory[22539] = 3'b110;
        rom_memory[22540] = 3'b111;
        rom_memory[22541] = 3'b111;
        rom_memory[22542] = 3'b111;
        rom_memory[22543] = 3'b111;
        rom_memory[22544] = 3'b111;
        rom_memory[22545] = 3'b110;
        rom_memory[22546] = 3'b110;
        rom_memory[22547] = 3'b110;
        rom_memory[22548] = 3'b111;
        rom_memory[22549] = 3'b110;
        rom_memory[22550] = 3'b111;
        rom_memory[22551] = 3'b111;
        rom_memory[22552] = 3'b111;
        rom_memory[22553] = 3'b110;
        rom_memory[22554] = 3'b110;
        rom_memory[22555] = 3'b110;
        rom_memory[22556] = 3'b110;
        rom_memory[22557] = 3'b110;
        rom_memory[22558] = 3'b110;
        rom_memory[22559] = 3'b110;
        rom_memory[22560] = 3'b110;
        rom_memory[22561] = 3'b110;
        rom_memory[22562] = 3'b110;
        rom_memory[22563] = 3'b110;
        rom_memory[22564] = 3'b110;
        rom_memory[22565] = 3'b110;
        rom_memory[22566] = 3'b110;
        rom_memory[22567] = 3'b110;
        rom_memory[22568] = 3'b110;
        rom_memory[22569] = 3'b110;
        rom_memory[22570] = 3'b110;
        rom_memory[22571] = 3'b110;
        rom_memory[22572] = 3'b110;
        rom_memory[22573] = 3'b110;
        rom_memory[22574] = 3'b110;
        rom_memory[22575] = 3'b110;
        rom_memory[22576] = 3'b110;
        rom_memory[22577] = 3'b110;
        rom_memory[22578] = 3'b110;
        rom_memory[22579] = 3'b110;
        rom_memory[22580] = 3'b110;
        rom_memory[22581] = 3'b110;
        rom_memory[22582] = 3'b110;
        rom_memory[22583] = 3'b110;
        rom_memory[22584] = 3'b110;
        rom_memory[22585] = 3'b110;
        rom_memory[22586] = 3'b110;
        rom_memory[22587] = 3'b110;
        rom_memory[22588] = 3'b110;
        rom_memory[22589] = 3'b111;
        rom_memory[22590] = 3'b111;
        rom_memory[22591] = 3'b111;
        rom_memory[22592] = 3'b111;
        rom_memory[22593] = 3'b111;
        rom_memory[22594] = 3'b111;
        rom_memory[22595] = 3'b111;
        rom_memory[22596] = 3'b111;
        rom_memory[22597] = 3'b111;
        rom_memory[22598] = 3'b111;
        rom_memory[22599] = 3'b111;
        rom_memory[22600] = 3'b111;
        rom_memory[22601] = 3'b111;
        rom_memory[22602] = 3'b111;
        rom_memory[22603] = 3'b111;
        rom_memory[22604] = 3'b111;
        rom_memory[22605] = 3'b111;
        rom_memory[22606] = 3'b111;
        rom_memory[22607] = 3'b111;
        rom_memory[22608] = 3'b111;
        rom_memory[22609] = 3'b110;
        rom_memory[22610] = 3'b100;
        rom_memory[22611] = 3'b100;
        rom_memory[22612] = 3'b100;
        rom_memory[22613] = 3'b110;
        rom_memory[22614] = 3'b110;
        rom_memory[22615] = 3'b100;
        rom_memory[22616] = 3'b100;
        rom_memory[22617] = 3'b100;
        rom_memory[22618] = 3'b100;
        rom_memory[22619] = 3'b100;
        rom_memory[22620] = 3'b100;
        rom_memory[22621] = 3'b100;
        rom_memory[22622] = 3'b110;
        rom_memory[22623] = 3'b110;
        rom_memory[22624] = 3'b110;
        rom_memory[22625] = 3'b100;
        rom_memory[22626] = 3'b110;
        rom_memory[22627] = 3'b110;
        rom_memory[22628] = 3'b110;
        rom_memory[22629] = 3'b110;
        rom_memory[22630] = 3'b110;
        rom_memory[22631] = 3'b110;
        rom_memory[22632] = 3'b110;
        rom_memory[22633] = 3'b110;
        rom_memory[22634] = 3'b110;
        rom_memory[22635] = 3'b110;
        rom_memory[22636] = 3'b110;
        rom_memory[22637] = 3'b110;
        rom_memory[22638] = 3'b110;
        rom_memory[22639] = 3'b110;
        rom_memory[22640] = 3'b110;
        rom_memory[22641] = 3'b110;
        rom_memory[22642] = 3'b110;
        rom_memory[22643] = 3'b110;
        rom_memory[22644] = 3'b110;
        rom_memory[22645] = 3'b110;
        rom_memory[22646] = 3'b110;
        rom_memory[22647] = 3'b110;
        rom_memory[22648] = 3'b110;
        rom_memory[22649] = 3'b110;
        rom_memory[22650] = 3'b110;
        rom_memory[22651] = 3'b110;
        rom_memory[22652] = 3'b110;
        rom_memory[22653] = 3'b110;
        rom_memory[22654] = 3'b110;
        rom_memory[22655] = 3'b110;
        rom_memory[22656] = 3'b110;
        rom_memory[22657] = 3'b110;
        rom_memory[22658] = 3'b110;
        rom_memory[22659] = 3'b110;
        rom_memory[22660] = 3'b110;
        rom_memory[22661] = 3'b111;
        rom_memory[22662] = 3'b111;
        rom_memory[22663] = 3'b111;
        rom_memory[22664] = 3'b111;
        rom_memory[22665] = 3'b111;
        rom_memory[22666] = 3'b111;
        rom_memory[22667] = 3'b111;
        rom_memory[22668] = 3'b111;
        rom_memory[22669] = 3'b111;
        rom_memory[22670] = 3'b110;
        rom_memory[22671] = 3'b000;
        rom_memory[22672] = 3'b000;
        rom_memory[22673] = 3'b000;
        rom_memory[22674] = 3'b000;
        rom_memory[22675] = 3'b000;
        rom_memory[22676] = 3'b000;
        rom_memory[22677] = 3'b000;
        rom_memory[22678] = 3'b100;
        rom_memory[22679] = 3'b000;
        rom_memory[22680] = 3'b100;
        rom_memory[22681] = 3'b000;
        rom_memory[22682] = 3'b100;
        rom_memory[22683] = 3'b110;
        rom_memory[22684] = 3'b110;
        rom_memory[22685] = 3'b110;
        rom_memory[22686] = 3'b111;
        rom_memory[22687] = 3'b111;
        rom_memory[22688] = 3'b111;
        rom_memory[22689] = 3'b110;
        rom_memory[22690] = 3'b110;
        rom_memory[22691] = 3'b110;
        rom_memory[22692] = 3'b110;
        rom_memory[22693] = 3'b110;
        rom_memory[22694] = 3'b110;
        rom_memory[22695] = 3'b110;
        rom_memory[22696] = 3'b110;
        rom_memory[22697] = 3'b110;
        rom_memory[22698] = 3'b110;
        rom_memory[22699] = 3'b110;
        rom_memory[22700] = 3'b110;
        rom_memory[22701] = 3'b110;
        rom_memory[22702] = 3'b110;
        rom_memory[22703] = 3'b110;
        rom_memory[22704] = 3'b110;
        rom_memory[22705] = 3'b110;
        rom_memory[22706] = 3'b110;
        rom_memory[22707] = 3'b110;
        rom_memory[22708] = 3'b110;
        rom_memory[22709] = 3'b110;
        rom_memory[22710] = 3'b110;
        rom_memory[22711] = 3'b111;
        rom_memory[22712] = 3'b111;
        rom_memory[22713] = 3'b111;
        rom_memory[22714] = 3'b111;
        rom_memory[22715] = 3'b111;
        rom_memory[22716] = 3'b111;
        rom_memory[22717] = 3'b111;
        rom_memory[22718] = 3'b111;
        rom_memory[22719] = 3'b111;
        rom_memory[22720] = 3'b111;
        rom_memory[22721] = 3'b111;
        rom_memory[22722] = 3'b111;
        rom_memory[22723] = 3'b111;
        rom_memory[22724] = 3'b111;
        rom_memory[22725] = 3'b111;
        rom_memory[22726] = 3'b111;
        rom_memory[22727] = 3'b111;
        rom_memory[22728] = 3'b111;
        rom_memory[22729] = 3'b111;
        rom_memory[22730] = 3'b111;
        rom_memory[22731] = 3'b111;
        rom_memory[22732] = 3'b111;
        rom_memory[22733] = 3'b111;
        rom_memory[22734] = 3'b111;
        rom_memory[22735] = 3'b111;
        rom_memory[22736] = 3'b111;
        rom_memory[22737] = 3'b111;
        rom_memory[22738] = 3'b111;
        rom_memory[22739] = 3'b111;
        rom_memory[22740] = 3'b111;
        rom_memory[22741] = 3'b111;
        rom_memory[22742] = 3'b111;
        rom_memory[22743] = 3'b111;
        rom_memory[22744] = 3'b111;
        rom_memory[22745] = 3'b111;
        rom_memory[22746] = 3'b111;
        rom_memory[22747] = 3'b110;
        rom_memory[22748] = 3'b110;
        rom_memory[22749] = 3'b110;
        rom_memory[22750] = 3'b111;
        rom_memory[22751] = 3'b111;
        rom_memory[22752] = 3'b110;
        rom_memory[22753] = 3'b110;
        rom_memory[22754] = 3'b110;
        rom_memory[22755] = 3'b110;
        rom_memory[22756] = 3'b110;
        rom_memory[22757] = 3'b110;
        rom_memory[22758] = 3'b111;
        rom_memory[22759] = 3'b111;
        rom_memory[22760] = 3'b111;
        rom_memory[22761] = 3'b111;
        rom_memory[22762] = 3'b111;
        rom_memory[22763] = 3'b111;
        rom_memory[22764] = 3'b111;
        rom_memory[22765] = 3'b111;
        rom_memory[22766] = 3'b111;
        rom_memory[22767] = 3'b111;
        rom_memory[22768] = 3'b111;
        rom_memory[22769] = 3'b111;
        rom_memory[22770] = 3'b110;
        rom_memory[22771] = 3'b111;
        rom_memory[22772] = 3'b111;
        rom_memory[22773] = 3'b111;
        rom_memory[22774] = 3'b110;
        rom_memory[22775] = 3'b111;
        rom_memory[22776] = 3'b110;
        rom_memory[22777] = 3'b110;
        rom_memory[22778] = 3'b111;
        rom_memory[22779] = 3'b111;
        rom_memory[22780] = 3'b111;
        rom_memory[22781] = 3'b111;
        rom_memory[22782] = 3'b111;
        rom_memory[22783] = 3'b111;
        rom_memory[22784] = 3'b111;
        rom_memory[22785] = 3'b110;
        rom_memory[22786] = 3'b110;
        rom_memory[22787] = 3'b110;
        rom_memory[22788] = 3'b111;
        rom_memory[22789] = 3'b111;
        rom_memory[22790] = 3'b111;
        rom_memory[22791] = 3'b110;
        rom_memory[22792] = 3'b110;
        rom_memory[22793] = 3'b111;
        rom_memory[22794] = 3'b110;
        rom_memory[22795] = 3'b111;
        rom_memory[22796] = 3'b111;
        rom_memory[22797] = 3'b111;
        rom_memory[22798] = 3'b110;
        rom_memory[22799] = 3'b110;
        rom_memory[22800] = 3'b110;
        rom_memory[22801] = 3'b110;
        rom_memory[22802] = 3'b110;
        rom_memory[22803] = 3'b110;
        rom_memory[22804] = 3'b110;
        rom_memory[22805] = 3'b110;
        rom_memory[22806] = 3'b110;
        rom_memory[22807] = 3'b110;
        rom_memory[22808] = 3'b110;
        rom_memory[22809] = 3'b110;
        rom_memory[22810] = 3'b110;
        rom_memory[22811] = 3'b110;
        rom_memory[22812] = 3'b110;
        rom_memory[22813] = 3'b110;
        rom_memory[22814] = 3'b110;
        rom_memory[22815] = 3'b110;
        rom_memory[22816] = 3'b110;
        rom_memory[22817] = 3'b110;
        rom_memory[22818] = 3'b110;
        rom_memory[22819] = 3'b110;
        rom_memory[22820] = 3'b110;
        rom_memory[22821] = 3'b110;
        rom_memory[22822] = 3'b110;
        rom_memory[22823] = 3'b110;
        rom_memory[22824] = 3'b110;
        rom_memory[22825] = 3'b110;
        rom_memory[22826] = 3'b110;
        rom_memory[22827] = 3'b110;
        rom_memory[22828] = 3'b110;
        rom_memory[22829] = 3'b111;
        rom_memory[22830] = 3'b111;
        rom_memory[22831] = 3'b111;
        rom_memory[22832] = 3'b111;
        rom_memory[22833] = 3'b111;
        rom_memory[22834] = 3'b111;
        rom_memory[22835] = 3'b111;
        rom_memory[22836] = 3'b111;
        rom_memory[22837] = 3'b111;
        rom_memory[22838] = 3'b111;
        rom_memory[22839] = 3'b111;
        rom_memory[22840] = 3'b111;
        rom_memory[22841] = 3'b111;
        rom_memory[22842] = 3'b111;
        rom_memory[22843] = 3'b111;
        rom_memory[22844] = 3'b111;
        rom_memory[22845] = 3'b111;
        rom_memory[22846] = 3'b111;
        rom_memory[22847] = 3'b111;
        rom_memory[22848] = 3'b111;
        rom_memory[22849] = 3'b110;
        rom_memory[22850] = 3'b100;
        rom_memory[22851] = 3'b100;
        rom_memory[22852] = 3'b100;
        rom_memory[22853] = 3'b110;
        rom_memory[22854] = 3'b110;
        rom_memory[22855] = 3'b100;
        rom_memory[22856] = 3'b100;
        rom_memory[22857] = 3'b100;
        rom_memory[22858] = 3'b100;
        rom_memory[22859] = 3'b100;
        rom_memory[22860] = 3'b100;
        rom_memory[22861] = 3'b100;
        rom_memory[22862] = 3'b100;
        rom_memory[22863] = 3'b110;
        rom_memory[22864] = 3'b110;
        rom_memory[22865] = 3'b110;
        rom_memory[22866] = 3'b110;
        rom_memory[22867] = 3'b110;
        rom_memory[22868] = 3'b110;
        rom_memory[22869] = 3'b110;
        rom_memory[22870] = 3'b110;
        rom_memory[22871] = 3'b110;
        rom_memory[22872] = 3'b110;
        rom_memory[22873] = 3'b110;
        rom_memory[22874] = 3'b110;
        rom_memory[22875] = 3'b110;
        rom_memory[22876] = 3'b110;
        rom_memory[22877] = 3'b110;
        rom_memory[22878] = 3'b110;
        rom_memory[22879] = 3'b110;
        rom_memory[22880] = 3'b110;
        rom_memory[22881] = 3'b110;
        rom_memory[22882] = 3'b110;
        rom_memory[22883] = 3'b110;
        rom_memory[22884] = 3'b110;
        rom_memory[22885] = 3'b110;
        rom_memory[22886] = 3'b110;
        rom_memory[22887] = 3'b110;
        rom_memory[22888] = 3'b110;
        rom_memory[22889] = 3'b110;
        rom_memory[22890] = 3'b110;
        rom_memory[22891] = 3'b110;
        rom_memory[22892] = 3'b110;
        rom_memory[22893] = 3'b110;
        rom_memory[22894] = 3'b110;
        rom_memory[22895] = 3'b110;
        rom_memory[22896] = 3'b110;
        rom_memory[22897] = 3'b110;
        rom_memory[22898] = 3'b110;
        rom_memory[22899] = 3'b110;
        rom_memory[22900] = 3'b110;
        rom_memory[22901] = 3'b110;
        rom_memory[22902] = 3'b111;
        rom_memory[22903] = 3'b111;
        rom_memory[22904] = 3'b111;
        rom_memory[22905] = 3'b111;
        rom_memory[22906] = 3'b111;
        rom_memory[22907] = 3'b111;
        rom_memory[22908] = 3'b111;
        rom_memory[22909] = 3'b111;
        rom_memory[22910] = 3'b111;
        rom_memory[22911] = 3'b111;
        rom_memory[22912] = 3'b100;
        rom_memory[22913] = 3'b000;
        rom_memory[22914] = 3'b000;
        rom_memory[22915] = 3'b000;
        rom_memory[22916] = 3'b000;
        rom_memory[22917] = 3'b000;
        rom_memory[22918] = 3'b000;
        rom_memory[22919] = 3'b100;
        rom_memory[22920] = 3'b000;
        rom_memory[22921] = 3'b100;
        rom_memory[22922] = 3'b000;
        rom_memory[22923] = 3'b100;
        rom_memory[22924] = 3'b110;
        rom_memory[22925] = 3'b110;
        rom_memory[22926] = 3'b111;
        rom_memory[22927] = 3'b111;
        rom_memory[22928] = 3'b111;
        rom_memory[22929] = 3'b111;
        rom_memory[22930] = 3'b110;
        rom_memory[22931] = 3'b110;
        rom_memory[22932] = 3'b110;
        rom_memory[22933] = 3'b110;
        rom_memory[22934] = 3'b110;
        rom_memory[22935] = 3'b110;
        rom_memory[22936] = 3'b110;
        rom_memory[22937] = 3'b110;
        rom_memory[22938] = 3'b110;
        rom_memory[22939] = 3'b110;
        rom_memory[22940] = 3'b110;
        rom_memory[22941] = 3'b110;
        rom_memory[22942] = 3'b110;
        rom_memory[22943] = 3'b110;
        rom_memory[22944] = 3'b110;
        rom_memory[22945] = 3'b110;
        rom_memory[22946] = 3'b110;
        rom_memory[22947] = 3'b111;
        rom_memory[22948] = 3'b110;
        rom_memory[22949] = 3'b110;
        rom_memory[22950] = 3'b110;
        rom_memory[22951] = 3'b110;
        rom_memory[22952] = 3'b110;
        rom_memory[22953] = 3'b111;
        rom_memory[22954] = 3'b111;
        rom_memory[22955] = 3'b111;
        rom_memory[22956] = 3'b111;
        rom_memory[22957] = 3'b111;
        rom_memory[22958] = 3'b111;
        rom_memory[22959] = 3'b111;
        rom_memory[22960] = 3'b111;
        rom_memory[22961] = 3'b111;
        rom_memory[22962] = 3'b110;
        rom_memory[22963] = 3'b111;
        rom_memory[22964] = 3'b111;
        rom_memory[22965] = 3'b111;
        rom_memory[22966] = 3'b111;
        rom_memory[22967] = 3'b111;
        rom_memory[22968] = 3'b111;
        rom_memory[22969] = 3'b111;
        rom_memory[22970] = 3'b111;
        rom_memory[22971] = 3'b111;
        rom_memory[22972] = 3'b111;
        rom_memory[22973] = 3'b111;
        rom_memory[22974] = 3'b111;
        rom_memory[22975] = 3'b111;
        rom_memory[22976] = 3'b111;
        rom_memory[22977] = 3'b111;
        rom_memory[22978] = 3'b111;
        rom_memory[22979] = 3'b111;
        rom_memory[22980] = 3'b111;
        rom_memory[22981] = 3'b111;
        rom_memory[22982] = 3'b111;
        rom_memory[22983] = 3'b111;
        rom_memory[22984] = 3'b111;
        rom_memory[22985] = 3'b111;
        rom_memory[22986] = 3'b111;
        rom_memory[22987] = 3'b111;
        rom_memory[22988] = 3'b111;
        rom_memory[22989] = 3'b111;
        rom_memory[22990] = 3'b111;
        rom_memory[22991] = 3'b111;
        rom_memory[22992] = 3'b111;
        rom_memory[22993] = 3'b111;
        rom_memory[22994] = 3'b110;
        rom_memory[22995] = 3'b110;
        rom_memory[22996] = 3'b111;
        rom_memory[22997] = 3'b111;
        rom_memory[22998] = 3'b111;
        rom_memory[22999] = 3'b111;
        rom_memory[23000] = 3'b111;
        rom_memory[23001] = 3'b111;
        rom_memory[23002] = 3'b111;
        rom_memory[23003] = 3'b111;
        rom_memory[23004] = 3'b111;
        rom_memory[23005] = 3'b111;
        rom_memory[23006] = 3'b111;
        rom_memory[23007] = 3'b111;
        rom_memory[23008] = 3'b111;
        rom_memory[23009] = 3'b111;
        rom_memory[23010] = 3'b111;
        rom_memory[23011] = 3'b111;
        rom_memory[23012] = 3'b111;
        rom_memory[23013] = 3'b111;
        rom_memory[23014] = 3'b111;
        rom_memory[23015] = 3'b111;
        rom_memory[23016] = 3'b111;
        rom_memory[23017] = 3'b111;
        rom_memory[23018] = 3'b111;
        rom_memory[23019] = 3'b111;
        rom_memory[23020] = 3'b111;
        rom_memory[23021] = 3'b111;
        rom_memory[23022] = 3'b111;
        rom_memory[23023] = 3'b111;
        rom_memory[23024] = 3'b111;
        rom_memory[23025] = 3'b111;
        rom_memory[23026] = 3'b111;
        rom_memory[23027] = 3'b111;
        rom_memory[23028] = 3'b111;
        rom_memory[23029] = 3'b110;
        rom_memory[23030] = 3'b111;
        rom_memory[23031] = 3'b111;
        rom_memory[23032] = 3'b111;
        rom_memory[23033] = 3'b111;
        rom_memory[23034] = 3'b110;
        rom_memory[23035] = 3'b111;
        rom_memory[23036] = 3'b111;
        rom_memory[23037] = 3'b111;
        rom_memory[23038] = 3'b110;
        rom_memory[23039] = 3'b110;
        rom_memory[23040] = 3'b110;
        rom_memory[23041] = 3'b110;
        rom_memory[23042] = 3'b110;
        rom_memory[23043] = 3'b110;
        rom_memory[23044] = 3'b110;
        rom_memory[23045] = 3'b110;
        rom_memory[23046] = 3'b110;
        rom_memory[23047] = 3'b110;
        rom_memory[23048] = 3'b110;
        rom_memory[23049] = 3'b110;
        rom_memory[23050] = 3'b110;
        rom_memory[23051] = 3'b110;
        rom_memory[23052] = 3'b110;
        rom_memory[23053] = 3'b110;
        rom_memory[23054] = 3'b110;
        rom_memory[23055] = 3'b110;
        rom_memory[23056] = 3'b110;
        rom_memory[23057] = 3'b110;
        rom_memory[23058] = 3'b110;
        rom_memory[23059] = 3'b110;
        rom_memory[23060] = 3'b110;
        rom_memory[23061] = 3'b110;
        rom_memory[23062] = 3'b110;
        rom_memory[23063] = 3'b110;
        rom_memory[23064] = 3'b110;
        rom_memory[23065] = 3'b110;
        rom_memory[23066] = 3'b110;
        rom_memory[23067] = 3'b110;
        rom_memory[23068] = 3'b111;
        rom_memory[23069] = 3'b111;
        rom_memory[23070] = 3'b111;
        rom_memory[23071] = 3'b111;
        rom_memory[23072] = 3'b111;
        rom_memory[23073] = 3'b111;
        rom_memory[23074] = 3'b111;
        rom_memory[23075] = 3'b111;
        rom_memory[23076] = 3'b111;
        rom_memory[23077] = 3'b111;
        rom_memory[23078] = 3'b111;
        rom_memory[23079] = 3'b111;
        rom_memory[23080] = 3'b111;
        rom_memory[23081] = 3'b111;
        rom_memory[23082] = 3'b111;
        rom_memory[23083] = 3'b111;
        rom_memory[23084] = 3'b111;
        rom_memory[23085] = 3'b111;
        rom_memory[23086] = 3'b111;
        rom_memory[23087] = 3'b111;
        rom_memory[23088] = 3'b111;
        rom_memory[23089] = 3'b111;
        rom_memory[23090] = 3'b100;
        rom_memory[23091] = 3'b100;
        rom_memory[23092] = 3'b100;
        rom_memory[23093] = 3'b100;
        rom_memory[23094] = 3'b110;
        rom_memory[23095] = 3'b100;
        rom_memory[23096] = 3'b100;
        rom_memory[23097] = 3'b100;
        rom_memory[23098] = 3'b100;
        rom_memory[23099] = 3'b100;
        rom_memory[23100] = 3'b100;
        rom_memory[23101] = 3'b100;
        rom_memory[23102] = 3'b100;
        rom_memory[23103] = 3'b110;
        rom_memory[23104] = 3'b110;
        rom_memory[23105] = 3'b110;
        rom_memory[23106] = 3'b110;
        rom_memory[23107] = 3'b110;
        rom_memory[23108] = 3'b110;
        rom_memory[23109] = 3'b110;
        rom_memory[23110] = 3'b110;
        rom_memory[23111] = 3'b110;
        rom_memory[23112] = 3'b110;
        rom_memory[23113] = 3'b110;
        rom_memory[23114] = 3'b110;
        rom_memory[23115] = 3'b110;
        rom_memory[23116] = 3'b110;
        rom_memory[23117] = 3'b110;
        rom_memory[23118] = 3'b110;
        rom_memory[23119] = 3'b110;
        rom_memory[23120] = 3'b110;
        rom_memory[23121] = 3'b110;
        rom_memory[23122] = 3'b110;
        rom_memory[23123] = 3'b110;
        rom_memory[23124] = 3'b110;
        rom_memory[23125] = 3'b110;
        rom_memory[23126] = 3'b110;
        rom_memory[23127] = 3'b110;
        rom_memory[23128] = 3'b110;
        rom_memory[23129] = 3'b110;
        rom_memory[23130] = 3'b110;
        rom_memory[23131] = 3'b110;
        rom_memory[23132] = 3'b110;
        rom_memory[23133] = 3'b110;
        rom_memory[23134] = 3'b110;
        rom_memory[23135] = 3'b110;
        rom_memory[23136] = 3'b110;
        rom_memory[23137] = 3'b110;
        rom_memory[23138] = 3'b110;
        rom_memory[23139] = 3'b110;
        rom_memory[23140] = 3'b110;
        rom_memory[23141] = 3'b110;
        rom_memory[23142] = 3'b110;
        rom_memory[23143] = 3'b111;
        rom_memory[23144] = 3'b111;
        rom_memory[23145] = 3'b111;
        rom_memory[23146] = 3'b111;
        rom_memory[23147] = 3'b111;
        rom_memory[23148] = 3'b111;
        rom_memory[23149] = 3'b111;
        rom_memory[23150] = 3'b111;
        rom_memory[23151] = 3'b111;
        rom_memory[23152] = 3'b111;
        rom_memory[23153] = 3'b111;
        rom_memory[23154] = 3'b000;
        rom_memory[23155] = 3'b000;
        rom_memory[23156] = 3'b000;
        rom_memory[23157] = 3'b000;
        rom_memory[23158] = 3'b000;
        rom_memory[23159] = 3'b000;
        rom_memory[23160] = 3'b100;
        rom_memory[23161] = 3'b000;
        rom_memory[23162] = 3'b100;
        rom_memory[23163] = 3'b000;
        rom_memory[23164] = 3'b100;
        rom_memory[23165] = 3'b110;
        rom_memory[23166] = 3'b111;
        rom_memory[23167] = 3'b111;
        rom_memory[23168] = 3'b111;
        rom_memory[23169] = 3'b111;
        rom_memory[23170] = 3'b110;
        rom_memory[23171] = 3'b110;
        rom_memory[23172] = 3'b110;
        rom_memory[23173] = 3'b110;
        rom_memory[23174] = 3'b110;
        rom_memory[23175] = 3'b110;
        rom_memory[23176] = 3'b110;
        rom_memory[23177] = 3'b110;
        rom_memory[23178] = 3'b110;
        rom_memory[23179] = 3'b110;
        rom_memory[23180] = 3'b110;
        rom_memory[23181] = 3'b110;
        rom_memory[23182] = 3'b110;
        rom_memory[23183] = 3'b110;
        rom_memory[23184] = 3'b110;
        rom_memory[23185] = 3'b110;
        rom_memory[23186] = 3'b110;
        rom_memory[23187] = 3'b110;
        rom_memory[23188] = 3'b110;
        rom_memory[23189] = 3'b110;
        rom_memory[23190] = 3'b110;
        rom_memory[23191] = 3'b110;
        rom_memory[23192] = 3'b110;
        rom_memory[23193] = 3'b111;
        rom_memory[23194] = 3'b111;
        rom_memory[23195] = 3'b111;
        rom_memory[23196] = 3'b111;
        rom_memory[23197] = 3'b110;
        rom_memory[23198] = 3'b110;
        rom_memory[23199] = 3'b111;
        rom_memory[23200] = 3'b110;
        rom_memory[23201] = 3'b111;
        rom_memory[23202] = 3'b111;
        rom_memory[23203] = 3'b111;
        rom_memory[23204] = 3'b111;
        rom_memory[23205] = 3'b111;
        rom_memory[23206] = 3'b111;
        rom_memory[23207] = 3'b111;
        rom_memory[23208] = 3'b111;
        rom_memory[23209] = 3'b111;
        rom_memory[23210] = 3'b111;
        rom_memory[23211] = 3'b111;
        rom_memory[23212] = 3'b111;
        rom_memory[23213] = 3'b111;
        rom_memory[23214] = 3'b111;
        rom_memory[23215] = 3'b111;
        rom_memory[23216] = 3'b111;
        rom_memory[23217] = 3'b111;
        rom_memory[23218] = 3'b111;
        rom_memory[23219] = 3'b111;
        rom_memory[23220] = 3'b111;
        rom_memory[23221] = 3'b111;
        rom_memory[23222] = 3'b111;
        rom_memory[23223] = 3'b111;
        rom_memory[23224] = 3'b111;
        rom_memory[23225] = 3'b111;
        rom_memory[23226] = 3'b111;
        rom_memory[23227] = 3'b111;
        rom_memory[23228] = 3'b111;
        rom_memory[23229] = 3'b111;
        rom_memory[23230] = 3'b111;
        rom_memory[23231] = 3'b111;
        rom_memory[23232] = 3'b111;
        rom_memory[23233] = 3'b111;
        rom_memory[23234] = 3'b111;
        rom_memory[23235] = 3'b111;
        rom_memory[23236] = 3'b111;
        rom_memory[23237] = 3'b111;
        rom_memory[23238] = 3'b111;
        rom_memory[23239] = 3'b111;
        rom_memory[23240] = 3'b111;
        rom_memory[23241] = 3'b111;
        rom_memory[23242] = 3'b111;
        rom_memory[23243] = 3'b111;
        rom_memory[23244] = 3'b111;
        rom_memory[23245] = 3'b111;
        rom_memory[23246] = 3'b111;
        rom_memory[23247] = 3'b111;
        rom_memory[23248] = 3'b111;
        rom_memory[23249] = 3'b111;
        rom_memory[23250] = 3'b111;
        rom_memory[23251] = 3'b111;
        rom_memory[23252] = 3'b111;
        rom_memory[23253] = 3'b111;
        rom_memory[23254] = 3'b111;
        rom_memory[23255] = 3'b111;
        rom_memory[23256] = 3'b111;
        rom_memory[23257] = 3'b111;
        rom_memory[23258] = 3'b111;
        rom_memory[23259] = 3'b111;
        rom_memory[23260] = 3'b111;
        rom_memory[23261] = 3'b111;
        rom_memory[23262] = 3'b111;
        rom_memory[23263] = 3'b111;
        rom_memory[23264] = 3'b111;
        rom_memory[23265] = 3'b111;
        rom_memory[23266] = 3'b111;
        rom_memory[23267] = 3'b111;
        rom_memory[23268] = 3'b111;
        rom_memory[23269] = 3'b111;
        rom_memory[23270] = 3'b111;
        rom_memory[23271] = 3'b111;
        rom_memory[23272] = 3'b111;
        rom_memory[23273] = 3'b111;
        rom_memory[23274] = 3'b111;
        rom_memory[23275] = 3'b111;
        rom_memory[23276] = 3'b111;
        rom_memory[23277] = 3'b111;
        rom_memory[23278] = 3'b111;
        rom_memory[23279] = 3'b111;
        rom_memory[23280] = 3'b110;
        rom_memory[23281] = 3'b110;
        rom_memory[23282] = 3'b110;
        rom_memory[23283] = 3'b110;
        rom_memory[23284] = 3'b110;
        rom_memory[23285] = 3'b110;
        rom_memory[23286] = 3'b110;
        rom_memory[23287] = 3'b110;
        rom_memory[23288] = 3'b110;
        rom_memory[23289] = 3'b110;
        rom_memory[23290] = 3'b110;
        rom_memory[23291] = 3'b110;
        rom_memory[23292] = 3'b110;
        rom_memory[23293] = 3'b110;
        rom_memory[23294] = 3'b110;
        rom_memory[23295] = 3'b110;
        rom_memory[23296] = 3'b110;
        rom_memory[23297] = 3'b110;
        rom_memory[23298] = 3'b110;
        rom_memory[23299] = 3'b110;
        rom_memory[23300] = 3'b110;
        rom_memory[23301] = 3'b110;
        rom_memory[23302] = 3'b110;
        rom_memory[23303] = 3'b110;
        rom_memory[23304] = 3'b110;
        rom_memory[23305] = 3'b110;
        rom_memory[23306] = 3'b110;
        rom_memory[23307] = 3'b110;
        rom_memory[23308] = 3'b111;
        rom_memory[23309] = 3'b111;
        rom_memory[23310] = 3'b111;
        rom_memory[23311] = 3'b111;
        rom_memory[23312] = 3'b111;
        rom_memory[23313] = 3'b111;
        rom_memory[23314] = 3'b111;
        rom_memory[23315] = 3'b111;
        rom_memory[23316] = 3'b111;
        rom_memory[23317] = 3'b111;
        rom_memory[23318] = 3'b111;
        rom_memory[23319] = 3'b111;
        rom_memory[23320] = 3'b111;
        rom_memory[23321] = 3'b111;
        rom_memory[23322] = 3'b111;
        rom_memory[23323] = 3'b111;
        rom_memory[23324] = 3'b111;
        rom_memory[23325] = 3'b111;
        rom_memory[23326] = 3'b111;
        rom_memory[23327] = 3'b111;
        rom_memory[23328] = 3'b111;
        rom_memory[23329] = 3'b111;
        rom_memory[23330] = 3'b110;
        rom_memory[23331] = 3'b100;
        rom_memory[23332] = 3'b100;
        rom_memory[23333] = 3'b100;
        rom_memory[23334] = 3'b100;
        rom_memory[23335] = 3'b100;
        rom_memory[23336] = 3'b100;
        rom_memory[23337] = 3'b100;
        rom_memory[23338] = 3'b100;
        rom_memory[23339] = 3'b100;
        rom_memory[23340] = 3'b100;
        rom_memory[23341] = 3'b100;
        rom_memory[23342] = 3'b110;
        rom_memory[23343] = 3'b110;
        rom_memory[23344] = 3'b110;
        rom_memory[23345] = 3'b110;
        rom_memory[23346] = 3'b110;
        rom_memory[23347] = 3'b110;
        rom_memory[23348] = 3'b110;
        rom_memory[23349] = 3'b110;
        rom_memory[23350] = 3'b110;
        rom_memory[23351] = 3'b110;
        rom_memory[23352] = 3'b110;
        rom_memory[23353] = 3'b110;
        rom_memory[23354] = 3'b110;
        rom_memory[23355] = 3'b110;
        rom_memory[23356] = 3'b110;
        rom_memory[23357] = 3'b110;
        rom_memory[23358] = 3'b110;
        rom_memory[23359] = 3'b110;
        rom_memory[23360] = 3'b110;
        rom_memory[23361] = 3'b110;
        rom_memory[23362] = 3'b110;
        rom_memory[23363] = 3'b110;
        rom_memory[23364] = 3'b110;
        rom_memory[23365] = 3'b110;
        rom_memory[23366] = 3'b110;
        rom_memory[23367] = 3'b110;
        rom_memory[23368] = 3'b110;
        rom_memory[23369] = 3'b110;
        rom_memory[23370] = 3'b110;
        rom_memory[23371] = 3'b110;
        rom_memory[23372] = 3'b110;
        rom_memory[23373] = 3'b110;
        rom_memory[23374] = 3'b110;
        rom_memory[23375] = 3'b110;
        rom_memory[23376] = 3'b110;
        rom_memory[23377] = 3'b110;
        rom_memory[23378] = 3'b110;
        rom_memory[23379] = 3'b110;
        rom_memory[23380] = 3'b110;
        rom_memory[23381] = 3'b110;
        rom_memory[23382] = 3'b110;
        rom_memory[23383] = 3'b110;
        rom_memory[23384] = 3'b111;
        rom_memory[23385] = 3'b111;
        rom_memory[23386] = 3'b111;
        rom_memory[23387] = 3'b111;
        rom_memory[23388] = 3'b111;
        rom_memory[23389] = 3'b111;
        rom_memory[23390] = 3'b111;
        rom_memory[23391] = 3'b111;
        rom_memory[23392] = 3'b111;
        rom_memory[23393] = 3'b111;
        rom_memory[23394] = 3'b111;
        rom_memory[23395] = 3'b100;
        rom_memory[23396] = 3'b000;
        rom_memory[23397] = 3'b000;
        rom_memory[23398] = 3'b000;
        rom_memory[23399] = 3'b000;
        rom_memory[23400] = 3'b000;
        rom_memory[23401] = 3'b100;
        rom_memory[23402] = 3'b000;
        rom_memory[23403] = 3'b100;
        rom_memory[23404] = 3'b000;
        rom_memory[23405] = 3'b110;
        rom_memory[23406] = 3'b110;
        rom_memory[23407] = 3'b111;
        rom_memory[23408] = 3'b110;
        rom_memory[23409] = 3'b110;
        rom_memory[23410] = 3'b110;
        rom_memory[23411] = 3'b110;
        rom_memory[23412] = 3'b110;
        rom_memory[23413] = 3'b110;
        rom_memory[23414] = 3'b110;
        rom_memory[23415] = 3'b110;
        rom_memory[23416] = 3'b110;
        rom_memory[23417] = 3'b110;
        rom_memory[23418] = 3'b110;
        rom_memory[23419] = 3'b110;
        rom_memory[23420] = 3'b110;
        rom_memory[23421] = 3'b110;
        rom_memory[23422] = 3'b110;
        rom_memory[23423] = 3'b110;
        rom_memory[23424] = 3'b110;
        rom_memory[23425] = 3'b110;
        rom_memory[23426] = 3'b110;
        rom_memory[23427] = 3'b110;
        rom_memory[23428] = 3'b110;
        rom_memory[23429] = 3'b110;
        rom_memory[23430] = 3'b110;
        rom_memory[23431] = 3'b110;
        rom_memory[23432] = 3'b110;
        rom_memory[23433] = 3'b111;
        rom_memory[23434] = 3'b111;
        rom_memory[23435] = 3'b110;
        rom_memory[23436] = 3'b110;
        rom_memory[23437] = 3'b110;
        rom_memory[23438] = 3'b110;
        rom_memory[23439] = 3'b110;
        rom_memory[23440] = 3'b110;
        rom_memory[23441] = 3'b110;
        rom_memory[23442] = 3'b111;
        rom_memory[23443] = 3'b111;
        rom_memory[23444] = 3'b111;
        rom_memory[23445] = 3'b111;
        rom_memory[23446] = 3'b111;
        rom_memory[23447] = 3'b111;
        rom_memory[23448] = 3'b111;
        rom_memory[23449] = 3'b111;
        rom_memory[23450] = 3'b111;
        rom_memory[23451] = 3'b111;
        rom_memory[23452] = 3'b111;
        rom_memory[23453] = 3'b111;
        rom_memory[23454] = 3'b111;
        rom_memory[23455] = 3'b111;
        rom_memory[23456] = 3'b111;
        rom_memory[23457] = 3'b111;
        rom_memory[23458] = 3'b111;
        rom_memory[23459] = 3'b111;
        rom_memory[23460] = 3'b111;
        rom_memory[23461] = 3'b111;
        rom_memory[23462] = 3'b111;
        rom_memory[23463] = 3'b111;
        rom_memory[23464] = 3'b111;
        rom_memory[23465] = 3'b111;
        rom_memory[23466] = 3'b111;
        rom_memory[23467] = 3'b111;
        rom_memory[23468] = 3'b111;
        rom_memory[23469] = 3'b111;
        rom_memory[23470] = 3'b111;
        rom_memory[23471] = 3'b111;
        rom_memory[23472] = 3'b111;
        rom_memory[23473] = 3'b111;
        rom_memory[23474] = 3'b111;
        rom_memory[23475] = 3'b111;
        rom_memory[23476] = 3'b111;
        rom_memory[23477] = 3'b111;
        rom_memory[23478] = 3'b111;
        rom_memory[23479] = 3'b111;
        rom_memory[23480] = 3'b111;
        rom_memory[23481] = 3'b111;
        rom_memory[23482] = 3'b111;
        rom_memory[23483] = 3'b111;
        rom_memory[23484] = 3'b111;
        rom_memory[23485] = 3'b111;
        rom_memory[23486] = 3'b111;
        rom_memory[23487] = 3'b111;
        rom_memory[23488] = 3'b111;
        rom_memory[23489] = 3'b111;
        rom_memory[23490] = 3'b111;
        rom_memory[23491] = 3'b111;
        rom_memory[23492] = 3'b111;
        rom_memory[23493] = 3'b111;
        rom_memory[23494] = 3'b111;
        rom_memory[23495] = 3'b111;
        rom_memory[23496] = 3'b111;
        rom_memory[23497] = 3'b111;
        rom_memory[23498] = 3'b111;
        rom_memory[23499] = 3'b111;
        rom_memory[23500] = 3'b111;
        rom_memory[23501] = 3'b111;
        rom_memory[23502] = 3'b111;
        rom_memory[23503] = 3'b111;
        rom_memory[23504] = 3'b111;
        rom_memory[23505] = 3'b111;
        rom_memory[23506] = 3'b111;
        rom_memory[23507] = 3'b111;
        rom_memory[23508] = 3'b111;
        rom_memory[23509] = 3'b111;
        rom_memory[23510] = 3'b111;
        rom_memory[23511] = 3'b111;
        rom_memory[23512] = 3'b111;
        rom_memory[23513] = 3'b111;
        rom_memory[23514] = 3'b111;
        rom_memory[23515] = 3'b111;
        rom_memory[23516] = 3'b111;
        rom_memory[23517] = 3'b111;
        rom_memory[23518] = 3'b111;
        rom_memory[23519] = 3'b111;
        rom_memory[23520] = 3'b110;
        rom_memory[23521] = 3'b110;
        rom_memory[23522] = 3'b110;
        rom_memory[23523] = 3'b110;
        rom_memory[23524] = 3'b110;
        rom_memory[23525] = 3'b110;
        rom_memory[23526] = 3'b110;
        rom_memory[23527] = 3'b110;
        rom_memory[23528] = 3'b110;
        rom_memory[23529] = 3'b110;
        rom_memory[23530] = 3'b110;
        rom_memory[23531] = 3'b110;
        rom_memory[23532] = 3'b110;
        rom_memory[23533] = 3'b110;
        rom_memory[23534] = 3'b110;
        rom_memory[23535] = 3'b110;
        rom_memory[23536] = 3'b110;
        rom_memory[23537] = 3'b110;
        rom_memory[23538] = 3'b110;
        rom_memory[23539] = 3'b110;
        rom_memory[23540] = 3'b110;
        rom_memory[23541] = 3'b110;
        rom_memory[23542] = 3'b110;
        rom_memory[23543] = 3'b110;
        rom_memory[23544] = 3'b110;
        rom_memory[23545] = 3'b110;
        rom_memory[23546] = 3'b110;
        rom_memory[23547] = 3'b110;
        rom_memory[23548] = 3'b111;
        rom_memory[23549] = 3'b111;
        rom_memory[23550] = 3'b111;
        rom_memory[23551] = 3'b111;
        rom_memory[23552] = 3'b111;
        rom_memory[23553] = 3'b111;
        rom_memory[23554] = 3'b111;
        rom_memory[23555] = 3'b111;
        rom_memory[23556] = 3'b111;
        rom_memory[23557] = 3'b111;
        rom_memory[23558] = 3'b111;
        rom_memory[23559] = 3'b111;
        rom_memory[23560] = 3'b111;
        rom_memory[23561] = 3'b111;
        rom_memory[23562] = 3'b111;
        rom_memory[23563] = 3'b111;
        rom_memory[23564] = 3'b111;
        rom_memory[23565] = 3'b111;
        rom_memory[23566] = 3'b111;
        rom_memory[23567] = 3'b111;
        rom_memory[23568] = 3'b111;
        rom_memory[23569] = 3'b111;
        rom_memory[23570] = 3'b110;
        rom_memory[23571] = 3'b110;
        rom_memory[23572] = 3'b100;
        rom_memory[23573] = 3'b100;
        rom_memory[23574] = 3'b100;
        rom_memory[23575] = 3'b100;
        rom_memory[23576] = 3'b100;
        rom_memory[23577] = 3'b100;
        rom_memory[23578] = 3'b100;
        rom_memory[23579] = 3'b100;
        rom_memory[23580] = 3'b100;
        rom_memory[23581] = 3'b100;
        rom_memory[23582] = 3'b110;
        rom_memory[23583] = 3'b110;
        rom_memory[23584] = 3'b110;
        rom_memory[23585] = 3'b110;
        rom_memory[23586] = 3'b110;
        rom_memory[23587] = 3'b110;
        rom_memory[23588] = 3'b110;
        rom_memory[23589] = 3'b110;
        rom_memory[23590] = 3'b110;
        rom_memory[23591] = 3'b110;
        rom_memory[23592] = 3'b110;
        rom_memory[23593] = 3'b110;
        rom_memory[23594] = 3'b110;
        rom_memory[23595] = 3'b110;
        rom_memory[23596] = 3'b110;
        rom_memory[23597] = 3'b110;
        rom_memory[23598] = 3'b110;
        rom_memory[23599] = 3'b110;
        rom_memory[23600] = 3'b110;
        rom_memory[23601] = 3'b110;
        rom_memory[23602] = 3'b110;
        rom_memory[23603] = 3'b110;
        rom_memory[23604] = 3'b110;
        rom_memory[23605] = 3'b110;
        rom_memory[23606] = 3'b110;
        rom_memory[23607] = 3'b110;
        rom_memory[23608] = 3'b110;
        rom_memory[23609] = 3'b110;
        rom_memory[23610] = 3'b110;
        rom_memory[23611] = 3'b110;
        rom_memory[23612] = 3'b110;
        rom_memory[23613] = 3'b110;
        rom_memory[23614] = 3'b110;
        rom_memory[23615] = 3'b110;
        rom_memory[23616] = 3'b110;
        rom_memory[23617] = 3'b110;
        rom_memory[23618] = 3'b110;
        rom_memory[23619] = 3'b110;
        rom_memory[23620] = 3'b110;
        rom_memory[23621] = 3'b110;
        rom_memory[23622] = 3'b110;
        rom_memory[23623] = 3'b110;
        rom_memory[23624] = 3'b111;
        rom_memory[23625] = 3'b111;
        rom_memory[23626] = 3'b111;
        rom_memory[23627] = 3'b111;
        rom_memory[23628] = 3'b111;
        rom_memory[23629] = 3'b111;
        rom_memory[23630] = 3'b111;
        rom_memory[23631] = 3'b111;
        rom_memory[23632] = 3'b111;
        rom_memory[23633] = 3'b111;
        rom_memory[23634] = 3'b111;
        rom_memory[23635] = 3'b111;
        rom_memory[23636] = 3'b000;
        rom_memory[23637] = 3'b000;
        rom_memory[23638] = 3'b000;
        rom_memory[23639] = 3'b000;
        rom_memory[23640] = 3'b000;
        rom_memory[23641] = 3'b000;
        rom_memory[23642] = 3'b100;
        rom_memory[23643] = 3'b000;
        rom_memory[23644] = 3'b100;
        rom_memory[23645] = 3'b100;
        rom_memory[23646] = 3'b110;
        rom_memory[23647] = 3'b110;
        rom_memory[23648] = 3'b110;
        rom_memory[23649] = 3'b110;
        rom_memory[23650] = 3'b110;
        rom_memory[23651] = 3'b110;
        rom_memory[23652] = 3'b110;
        rom_memory[23653] = 3'b110;
        rom_memory[23654] = 3'b110;
        rom_memory[23655] = 3'b110;
        rom_memory[23656] = 3'b110;
        rom_memory[23657] = 3'b110;
        rom_memory[23658] = 3'b110;
        rom_memory[23659] = 3'b110;
        rom_memory[23660] = 3'b110;
        rom_memory[23661] = 3'b110;
        rom_memory[23662] = 3'b110;
        rom_memory[23663] = 3'b110;
        rom_memory[23664] = 3'b110;
        rom_memory[23665] = 3'b110;
        rom_memory[23666] = 3'b110;
        rom_memory[23667] = 3'b110;
        rom_memory[23668] = 3'b110;
        rom_memory[23669] = 3'b110;
        rom_memory[23670] = 3'b110;
        rom_memory[23671] = 3'b110;
        rom_memory[23672] = 3'b110;
        rom_memory[23673] = 3'b110;
        rom_memory[23674] = 3'b110;
        rom_memory[23675] = 3'b110;
        rom_memory[23676] = 3'b110;
        rom_memory[23677] = 3'b110;
        rom_memory[23678] = 3'b110;
        rom_memory[23679] = 3'b111;
        rom_memory[23680] = 3'b110;
        rom_memory[23681] = 3'b110;
        rom_memory[23682] = 3'b111;
        rom_memory[23683] = 3'b111;
        rom_memory[23684] = 3'b111;
        rom_memory[23685] = 3'b111;
        rom_memory[23686] = 3'b111;
        rom_memory[23687] = 3'b111;
        rom_memory[23688] = 3'b111;
        rom_memory[23689] = 3'b111;
        rom_memory[23690] = 3'b111;
        rom_memory[23691] = 3'b111;
        rom_memory[23692] = 3'b111;
        rom_memory[23693] = 3'b111;
        rom_memory[23694] = 3'b111;
        rom_memory[23695] = 3'b111;
        rom_memory[23696] = 3'b111;
        rom_memory[23697] = 3'b111;
        rom_memory[23698] = 3'b111;
        rom_memory[23699] = 3'b111;
        rom_memory[23700] = 3'b111;
        rom_memory[23701] = 3'b111;
        rom_memory[23702] = 3'b111;
        rom_memory[23703] = 3'b111;
        rom_memory[23704] = 3'b111;
        rom_memory[23705] = 3'b111;
        rom_memory[23706] = 3'b111;
        rom_memory[23707] = 3'b111;
        rom_memory[23708] = 3'b111;
        rom_memory[23709] = 3'b111;
        rom_memory[23710] = 3'b111;
        rom_memory[23711] = 3'b111;
        rom_memory[23712] = 3'b111;
        rom_memory[23713] = 3'b111;
        rom_memory[23714] = 3'b111;
        rom_memory[23715] = 3'b111;
        rom_memory[23716] = 3'b111;
        rom_memory[23717] = 3'b111;
        rom_memory[23718] = 3'b111;
        rom_memory[23719] = 3'b111;
        rom_memory[23720] = 3'b111;
        rom_memory[23721] = 3'b111;
        rom_memory[23722] = 3'b111;
        rom_memory[23723] = 3'b111;
        rom_memory[23724] = 3'b111;
        rom_memory[23725] = 3'b111;
        rom_memory[23726] = 3'b111;
        rom_memory[23727] = 3'b111;
        rom_memory[23728] = 3'b111;
        rom_memory[23729] = 3'b111;
        rom_memory[23730] = 3'b111;
        rom_memory[23731] = 3'b111;
        rom_memory[23732] = 3'b111;
        rom_memory[23733] = 3'b111;
        rom_memory[23734] = 3'b111;
        rom_memory[23735] = 3'b111;
        rom_memory[23736] = 3'b111;
        rom_memory[23737] = 3'b111;
        rom_memory[23738] = 3'b111;
        rom_memory[23739] = 3'b111;
        rom_memory[23740] = 3'b111;
        rom_memory[23741] = 3'b111;
        rom_memory[23742] = 3'b111;
        rom_memory[23743] = 3'b111;
        rom_memory[23744] = 3'b111;
        rom_memory[23745] = 3'b111;
        rom_memory[23746] = 3'b111;
        rom_memory[23747] = 3'b111;
        rom_memory[23748] = 3'b111;
        rom_memory[23749] = 3'b111;
        rom_memory[23750] = 3'b111;
        rom_memory[23751] = 3'b111;
        rom_memory[23752] = 3'b111;
        rom_memory[23753] = 3'b111;
        rom_memory[23754] = 3'b111;
        rom_memory[23755] = 3'b111;
        rom_memory[23756] = 3'b111;
        rom_memory[23757] = 3'b111;
        rom_memory[23758] = 3'b111;
        rom_memory[23759] = 3'b111;
        rom_memory[23760] = 3'b110;
        rom_memory[23761] = 3'b110;
        rom_memory[23762] = 3'b110;
        rom_memory[23763] = 3'b110;
        rom_memory[23764] = 3'b110;
        rom_memory[23765] = 3'b110;
        rom_memory[23766] = 3'b110;
        rom_memory[23767] = 3'b110;
        rom_memory[23768] = 3'b110;
        rom_memory[23769] = 3'b110;
        rom_memory[23770] = 3'b110;
        rom_memory[23771] = 3'b110;
        rom_memory[23772] = 3'b110;
        rom_memory[23773] = 3'b110;
        rom_memory[23774] = 3'b110;
        rom_memory[23775] = 3'b110;
        rom_memory[23776] = 3'b110;
        rom_memory[23777] = 3'b110;
        rom_memory[23778] = 3'b110;
        rom_memory[23779] = 3'b110;
        rom_memory[23780] = 3'b110;
        rom_memory[23781] = 3'b110;
        rom_memory[23782] = 3'b110;
        rom_memory[23783] = 3'b110;
        rom_memory[23784] = 3'b110;
        rom_memory[23785] = 3'b110;
        rom_memory[23786] = 3'b110;
        rom_memory[23787] = 3'b111;
        rom_memory[23788] = 3'b111;
        rom_memory[23789] = 3'b111;
        rom_memory[23790] = 3'b111;
        rom_memory[23791] = 3'b111;
        rom_memory[23792] = 3'b111;
        rom_memory[23793] = 3'b111;
        rom_memory[23794] = 3'b111;
        rom_memory[23795] = 3'b111;
        rom_memory[23796] = 3'b111;
        rom_memory[23797] = 3'b111;
        rom_memory[23798] = 3'b111;
        rom_memory[23799] = 3'b111;
        rom_memory[23800] = 3'b111;
        rom_memory[23801] = 3'b111;
        rom_memory[23802] = 3'b111;
        rom_memory[23803] = 3'b111;
        rom_memory[23804] = 3'b111;
        rom_memory[23805] = 3'b111;
        rom_memory[23806] = 3'b111;
        rom_memory[23807] = 3'b111;
        rom_memory[23808] = 3'b111;
        rom_memory[23809] = 3'b111;
        rom_memory[23810] = 3'b111;
        rom_memory[23811] = 3'b110;
        rom_memory[23812] = 3'b100;
        rom_memory[23813] = 3'b100;
        rom_memory[23814] = 3'b100;
        rom_memory[23815] = 3'b100;
        rom_memory[23816] = 3'b100;
        rom_memory[23817] = 3'b100;
        rom_memory[23818] = 3'b100;
        rom_memory[23819] = 3'b100;
        rom_memory[23820] = 3'b100;
        rom_memory[23821] = 3'b100;
        rom_memory[23822] = 3'b100;
        rom_memory[23823] = 3'b110;
        rom_memory[23824] = 3'b110;
        rom_memory[23825] = 3'b110;
        rom_memory[23826] = 3'b110;
        rom_memory[23827] = 3'b110;
        rom_memory[23828] = 3'b110;
        rom_memory[23829] = 3'b110;
        rom_memory[23830] = 3'b110;
        rom_memory[23831] = 3'b110;
        rom_memory[23832] = 3'b110;
        rom_memory[23833] = 3'b110;
        rom_memory[23834] = 3'b110;
        rom_memory[23835] = 3'b110;
        rom_memory[23836] = 3'b110;
        rom_memory[23837] = 3'b110;
        rom_memory[23838] = 3'b110;
        rom_memory[23839] = 3'b110;
        rom_memory[23840] = 3'b110;
        rom_memory[23841] = 3'b110;
        rom_memory[23842] = 3'b110;
        rom_memory[23843] = 3'b110;
        rom_memory[23844] = 3'b110;
        rom_memory[23845] = 3'b110;
        rom_memory[23846] = 3'b110;
        rom_memory[23847] = 3'b110;
        rom_memory[23848] = 3'b110;
        rom_memory[23849] = 3'b110;
        rom_memory[23850] = 3'b110;
        rom_memory[23851] = 3'b110;
        rom_memory[23852] = 3'b110;
        rom_memory[23853] = 3'b110;
        rom_memory[23854] = 3'b110;
        rom_memory[23855] = 3'b110;
        rom_memory[23856] = 3'b110;
        rom_memory[23857] = 3'b110;
        rom_memory[23858] = 3'b110;
        rom_memory[23859] = 3'b110;
        rom_memory[23860] = 3'b110;
        rom_memory[23861] = 3'b110;
        rom_memory[23862] = 3'b110;
        rom_memory[23863] = 3'b110;
        rom_memory[23864] = 3'b110;
        rom_memory[23865] = 3'b111;
        rom_memory[23866] = 3'b111;
        rom_memory[23867] = 3'b111;
        rom_memory[23868] = 3'b111;
        rom_memory[23869] = 3'b111;
        rom_memory[23870] = 3'b111;
        rom_memory[23871] = 3'b111;
        rom_memory[23872] = 3'b111;
        rom_memory[23873] = 3'b111;
        rom_memory[23874] = 3'b111;
        rom_memory[23875] = 3'b111;
        rom_memory[23876] = 3'b110;
        rom_memory[23877] = 3'b000;
        rom_memory[23878] = 3'b000;
        rom_memory[23879] = 3'b000;
        rom_memory[23880] = 3'b000;
        rom_memory[23881] = 3'b000;
        rom_memory[23882] = 3'b000;
        rom_memory[23883] = 3'b100;
        rom_memory[23884] = 3'b100;
        rom_memory[23885] = 3'b000;
        rom_memory[23886] = 3'b100;
        rom_memory[23887] = 3'b110;
        rom_memory[23888] = 3'b110;
        rom_memory[23889] = 3'b110;
        rom_memory[23890] = 3'b110;
        rom_memory[23891] = 3'b110;
        rom_memory[23892] = 3'b110;
        rom_memory[23893] = 3'b110;
        rom_memory[23894] = 3'b110;
        rom_memory[23895] = 3'b110;
        rom_memory[23896] = 3'b110;
        rom_memory[23897] = 3'b110;
        rom_memory[23898] = 3'b110;
        rom_memory[23899] = 3'b110;
        rom_memory[23900] = 3'b110;
        rom_memory[23901] = 3'b110;
        rom_memory[23902] = 3'b110;
        rom_memory[23903] = 3'b110;
        rom_memory[23904] = 3'b110;
        rom_memory[23905] = 3'b110;
        rom_memory[23906] = 3'b110;
        rom_memory[23907] = 3'b110;
        rom_memory[23908] = 3'b110;
        rom_memory[23909] = 3'b110;
        rom_memory[23910] = 3'b110;
        rom_memory[23911] = 3'b110;
        rom_memory[23912] = 3'b110;
        rom_memory[23913] = 3'b110;
        rom_memory[23914] = 3'b110;
        rom_memory[23915] = 3'b110;
        rom_memory[23916] = 3'b110;
        rom_memory[23917] = 3'b110;
        rom_memory[23918] = 3'b110;
        rom_memory[23919] = 3'b111;
        rom_memory[23920] = 3'b110;
        rom_memory[23921] = 3'b110;
        rom_memory[23922] = 3'b111;
        rom_memory[23923] = 3'b111;
        rom_memory[23924] = 3'b111;
        rom_memory[23925] = 3'b111;
        rom_memory[23926] = 3'b111;
        rom_memory[23927] = 3'b111;
        rom_memory[23928] = 3'b111;
        rom_memory[23929] = 3'b111;
        rom_memory[23930] = 3'b111;
        rom_memory[23931] = 3'b111;
        rom_memory[23932] = 3'b111;
        rom_memory[23933] = 3'b111;
        rom_memory[23934] = 3'b111;
        rom_memory[23935] = 3'b111;
        rom_memory[23936] = 3'b111;
        rom_memory[23937] = 3'b111;
        rom_memory[23938] = 3'b111;
        rom_memory[23939] = 3'b111;
        rom_memory[23940] = 3'b111;
        rom_memory[23941] = 3'b111;
        rom_memory[23942] = 3'b111;
        rom_memory[23943] = 3'b111;
        rom_memory[23944] = 3'b111;
        rom_memory[23945] = 3'b111;
        rom_memory[23946] = 3'b110;
        rom_memory[23947] = 3'b111;
        rom_memory[23948] = 3'b111;
        rom_memory[23949] = 3'b111;
        rom_memory[23950] = 3'b111;
        rom_memory[23951] = 3'b111;
        rom_memory[23952] = 3'b111;
        rom_memory[23953] = 3'b111;
        rom_memory[23954] = 3'b111;
        rom_memory[23955] = 3'b111;
        rom_memory[23956] = 3'b111;
        rom_memory[23957] = 3'b111;
        rom_memory[23958] = 3'b111;
        rom_memory[23959] = 3'b111;
        rom_memory[23960] = 3'b111;
        rom_memory[23961] = 3'b111;
        rom_memory[23962] = 3'b111;
        rom_memory[23963] = 3'b111;
        rom_memory[23964] = 3'b111;
        rom_memory[23965] = 3'b111;
        rom_memory[23966] = 3'b111;
        rom_memory[23967] = 3'b111;
        rom_memory[23968] = 3'b111;
        rom_memory[23969] = 3'b111;
        rom_memory[23970] = 3'b111;
        rom_memory[23971] = 3'b111;
        rom_memory[23972] = 3'b111;
        rom_memory[23973] = 3'b111;
        rom_memory[23974] = 3'b111;
        rom_memory[23975] = 3'b111;
        rom_memory[23976] = 3'b111;
        rom_memory[23977] = 3'b111;
        rom_memory[23978] = 3'b111;
        rom_memory[23979] = 3'b111;
        rom_memory[23980] = 3'b111;
        rom_memory[23981] = 3'b111;
        rom_memory[23982] = 3'b111;
        rom_memory[23983] = 3'b111;
        rom_memory[23984] = 3'b111;
        rom_memory[23985] = 3'b111;
        rom_memory[23986] = 3'b111;
        rom_memory[23987] = 3'b111;
        rom_memory[23988] = 3'b111;
        rom_memory[23989] = 3'b111;
        rom_memory[23990] = 3'b111;
        rom_memory[23991] = 3'b111;
        rom_memory[23992] = 3'b111;
        rom_memory[23993] = 3'b111;
        rom_memory[23994] = 3'b111;
        rom_memory[23995] = 3'b111;
        rom_memory[23996] = 3'b111;
        rom_memory[23997] = 3'b111;
        rom_memory[23998] = 3'b111;
        rom_memory[23999] = 3'b111;
        rom_memory[24000] = 3'b110;
        rom_memory[24001] = 3'b110;
        rom_memory[24002] = 3'b110;
        rom_memory[24003] = 3'b110;
        rom_memory[24004] = 3'b110;
        rom_memory[24005] = 3'b110;
        rom_memory[24006] = 3'b110;
        rom_memory[24007] = 3'b110;
        rom_memory[24008] = 3'b110;
        rom_memory[24009] = 3'b110;
        rom_memory[24010] = 3'b110;
        rom_memory[24011] = 3'b110;
        rom_memory[24012] = 3'b110;
        rom_memory[24013] = 3'b110;
        rom_memory[24014] = 3'b110;
        rom_memory[24015] = 3'b110;
        rom_memory[24016] = 3'b110;
        rom_memory[24017] = 3'b110;
        rom_memory[24018] = 3'b110;
        rom_memory[24019] = 3'b110;
        rom_memory[24020] = 3'b110;
        rom_memory[24021] = 3'b110;
        rom_memory[24022] = 3'b110;
        rom_memory[24023] = 3'b110;
        rom_memory[24024] = 3'b110;
        rom_memory[24025] = 3'b110;
        rom_memory[24026] = 3'b110;
        rom_memory[24027] = 3'b111;
        rom_memory[24028] = 3'b111;
        rom_memory[24029] = 3'b111;
        rom_memory[24030] = 3'b111;
        rom_memory[24031] = 3'b111;
        rom_memory[24032] = 3'b111;
        rom_memory[24033] = 3'b111;
        rom_memory[24034] = 3'b111;
        rom_memory[24035] = 3'b111;
        rom_memory[24036] = 3'b111;
        rom_memory[24037] = 3'b111;
        rom_memory[24038] = 3'b111;
        rom_memory[24039] = 3'b111;
        rom_memory[24040] = 3'b111;
        rom_memory[24041] = 3'b111;
        rom_memory[24042] = 3'b111;
        rom_memory[24043] = 3'b111;
        rom_memory[24044] = 3'b111;
        rom_memory[24045] = 3'b111;
        rom_memory[24046] = 3'b111;
        rom_memory[24047] = 3'b111;
        rom_memory[24048] = 3'b111;
        rom_memory[24049] = 3'b111;
        rom_memory[24050] = 3'b111;
        rom_memory[24051] = 3'b110;
        rom_memory[24052] = 3'b110;
        rom_memory[24053] = 3'b100;
        rom_memory[24054] = 3'b100;
        rom_memory[24055] = 3'b100;
        rom_memory[24056] = 3'b100;
        rom_memory[24057] = 3'b100;
        rom_memory[24058] = 3'b100;
        rom_memory[24059] = 3'b100;
        rom_memory[24060] = 3'b100;
        rom_memory[24061] = 3'b100;
        rom_memory[24062] = 3'b100;
        rom_memory[24063] = 3'b110;
        rom_memory[24064] = 3'b110;
        rom_memory[24065] = 3'b110;
        rom_memory[24066] = 3'b110;
        rom_memory[24067] = 3'b110;
        rom_memory[24068] = 3'b110;
        rom_memory[24069] = 3'b110;
        rom_memory[24070] = 3'b110;
        rom_memory[24071] = 3'b110;
        rom_memory[24072] = 3'b110;
        rom_memory[24073] = 3'b110;
        rom_memory[24074] = 3'b110;
        rom_memory[24075] = 3'b110;
        rom_memory[24076] = 3'b110;
        rom_memory[24077] = 3'b110;
        rom_memory[24078] = 3'b110;
        rom_memory[24079] = 3'b110;
        rom_memory[24080] = 3'b110;
        rom_memory[24081] = 3'b110;
        rom_memory[24082] = 3'b110;
        rom_memory[24083] = 3'b110;
        rom_memory[24084] = 3'b110;
        rom_memory[24085] = 3'b110;
        rom_memory[24086] = 3'b110;
        rom_memory[24087] = 3'b110;
        rom_memory[24088] = 3'b110;
        rom_memory[24089] = 3'b110;
        rom_memory[24090] = 3'b110;
        rom_memory[24091] = 3'b110;
        rom_memory[24092] = 3'b110;
        rom_memory[24093] = 3'b110;
        rom_memory[24094] = 3'b110;
        rom_memory[24095] = 3'b110;
        rom_memory[24096] = 3'b110;
        rom_memory[24097] = 3'b110;
        rom_memory[24098] = 3'b110;
        rom_memory[24099] = 3'b110;
        rom_memory[24100] = 3'b110;
        rom_memory[24101] = 3'b110;
        rom_memory[24102] = 3'b110;
        rom_memory[24103] = 3'b110;
        rom_memory[24104] = 3'b110;
        rom_memory[24105] = 3'b111;
        rom_memory[24106] = 3'b111;
        rom_memory[24107] = 3'b111;
        rom_memory[24108] = 3'b111;
        rom_memory[24109] = 3'b111;
        rom_memory[24110] = 3'b111;
        rom_memory[24111] = 3'b111;
        rom_memory[24112] = 3'b111;
        rom_memory[24113] = 3'b111;
        rom_memory[24114] = 3'b111;
        rom_memory[24115] = 3'b111;
        rom_memory[24116] = 3'b111;
        rom_memory[24117] = 3'b110;
        rom_memory[24118] = 3'b000;
        rom_memory[24119] = 3'b000;
        rom_memory[24120] = 3'b000;
        rom_memory[24121] = 3'b000;
        rom_memory[24122] = 3'b000;
        rom_memory[24123] = 3'b000;
        rom_memory[24124] = 3'b000;
        rom_memory[24125] = 3'b000;
        rom_memory[24126] = 3'b000;
        rom_memory[24127] = 3'b110;
        rom_memory[24128] = 3'b111;
        rom_memory[24129] = 3'b110;
        rom_memory[24130] = 3'b110;
        rom_memory[24131] = 3'b110;
        rom_memory[24132] = 3'b110;
        rom_memory[24133] = 3'b110;
        rom_memory[24134] = 3'b110;
        rom_memory[24135] = 3'b110;
        rom_memory[24136] = 3'b110;
        rom_memory[24137] = 3'b110;
        rom_memory[24138] = 3'b110;
        rom_memory[24139] = 3'b110;
        rom_memory[24140] = 3'b110;
        rom_memory[24141] = 3'b110;
        rom_memory[24142] = 3'b110;
        rom_memory[24143] = 3'b110;
        rom_memory[24144] = 3'b110;
        rom_memory[24145] = 3'b110;
        rom_memory[24146] = 3'b110;
        rom_memory[24147] = 3'b110;
        rom_memory[24148] = 3'b110;
        rom_memory[24149] = 3'b110;
        rom_memory[24150] = 3'b110;
        rom_memory[24151] = 3'b110;
        rom_memory[24152] = 3'b110;
        rom_memory[24153] = 3'b110;
        rom_memory[24154] = 3'b110;
        rom_memory[24155] = 3'b110;
        rom_memory[24156] = 3'b110;
        rom_memory[24157] = 3'b110;
        rom_memory[24158] = 3'b110;
        rom_memory[24159] = 3'b110;
        rom_memory[24160] = 3'b110;
        rom_memory[24161] = 3'b110;
        rom_memory[24162] = 3'b111;
        rom_memory[24163] = 3'b110;
        rom_memory[24164] = 3'b111;
        rom_memory[24165] = 3'b111;
        rom_memory[24166] = 3'b111;
        rom_memory[24167] = 3'b111;
        rom_memory[24168] = 3'b111;
        rom_memory[24169] = 3'b111;
        rom_memory[24170] = 3'b111;
        rom_memory[24171] = 3'b111;
        rom_memory[24172] = 3'b111;
        rom_memory[24173] = 3'b111;
        rom_memory[24174] = 3'b111;
        rom_memory[24175] = 3'b111;
        rom_memory[24176] = 3'b111;
        rom_memory[24177] = 3'b111;
        rom_memory[24178] = 3'b111;
        rom_memory[24179] = 3'b111;
        rom_memory[24180] = 3'b111;
        rom_memory[24181] = 3'b111;
        rom_memory[24182] = 3'b111;
        rom_memory[24183] = 3'b111;
        rom_memory[24184] = 3'b111;
        rom_memory[24185] = 3'b111;
        rom_memory[24186] = 3'b110;
        rom_memory[24187] = 3'b110;
        rom_memory[24188] = 3'b111;
        rom_memory[24189] = 3'b111;
        rom_memory[24190] = 3'b111;
        rom_memory[24191] = 3'b111;
        rom_memory[24192] = 3'b111;
        rom_memory[24193] = 3'b111;
        rom_memory[24194] = 3'b111;
        rom_memory[24195] = 3'b111;
        rom_memory[24196] = 3'b111;
        rom_memory[24197] = 3'b111;
        rom_memory[24198] = 3'b111;
        rom_memory[24199] = 3'b111;
        rom_memory[24200] = 3'b111;
        rom_memory[24201] = 3'b111;
        rom_memory[24202] = 3'b111;
        rom_memory[24203] = 3'b111;
        rom_memory[24204] = 3'b111;
        rom_memory[24205] = 3'b111;
        rom_memory[24206] = 3'b111;
        rom_memory[24207] = 3'b111;
        rom_memory[24208] = 3'b111;
        rom_memory[24209] = 3'b111;
        rom_memory[24210] = 3'b111;
        rom_memory[24211] = 3'b111;
        rom_memory[24212] = 3'b111;
        rom_memory[24213] = 3'b111;
        rom_memory[24214] = 3'b111;
        rom_memory[24215] = 3'b111;
        rom_memory[24216] = 3'b111;
        rom_memory[24217] = 3'b111;
        rom_memory[24218] = 3'b111;
        rom_memory[24219] = 3'b111;
        rom_memory[24220] = 3'b111;
        rom_memory[24221] = 3'b111;
        rom_memory[24222] = 3'b111;
        rom_memory[24223] = 3'b111;
        rom_memory[24224] = 3'b111;
        rom_memory[24225] = 3'b111;
        rom_memory[24226] = 3'b111;
        rom_memory[24227] = 3'b111;
        rom_memory[24228] = 3'b111;
        rom_memory[24229] = 3'b111;
        rom_memory[24230] = 3'b111;
        rom_memory[24231] = 3'b111;
        rom_memory[24232] = 3'b111;
        rom_memory[24233] = 3'b111;
        rom_memory[24234] = 3'b111;
        rom_memory[24235] = 3'b111;
        rom_memory[24236] = 3'b111;
        rom_memory[24237] = 3'b111;
        rom_memory[24238] = 3'b111;
        rom_memory[24239] = 3'b111;
        rom_memory[24240] = 3'b110;
        rom_memory[24241] = 3'b110;
        rom_memory[24242] = 3'b110;
        rom_memory[24243] = 3'b110;
        rom_memory[24244] = 3'b110;
        rom_memory[24245] = 3'b110;
        rom_memory[24246] = 3'b110;
        rom_memory[24247] = 3'b110;
        rom_memory[24248] = 3'b110;
        rom_memory[24249] = 3'b110;
        rom_memory[24250] = 3'b110;
        rom_memory[24251] = 3'b110;
        rom_memory[24252] = 3'b110;
        rom_memory[24253] = 3'b110;
        rom_memory[24254] = 3'b110;
        rom_memory[24255] = 3'b110;
        rom_memory[24256] = 3'b110;
        rom_memory[24257] = 3'b110;
        rom_memory[24258] = 3'b110;
        rom_memory[24259] = 3'b110;
        rom_memory[24260] = 3'b110;
        rom_memory[24261] = 3'b110;
        rom_memory[24262] = 3'b110;
        rom_memory[24263] = 3'b110;
        rom_memory[24264] = 3'b110;
        rom_memory[24265] = 3'b110;
        rom_memory[24266] = 3'b110;
        rom_memory[24267] = 3'b110;
        rom_memory[24268] = 3'b111;
        rom_memory[24269] = 3'b111;
        rom_memory[24270] = 3'b111;
        rom_memory[24271] = 3'b111;
        rom_memory[24272] = 3'b111;
        rom_memory[24273] = 3'b111;
        rom_memory[24274] = 3'b111;
        rom_memory[24275] = 3'b111;
        rom_memory[24276] = 3'b111;
        rom_memory[24277] = 3'b111;
        rom_memory[24278] = 3'b111;
        rom_memory[24279] = 3'b111;
        rom_memory[24280] = 3'b111;
        rom_memory[24281] = 3'b111;
        rom_memory[24282] = 3'b111;
        rom_memory[24283] = 3'b111;
        rom_memory[24284] = 3'b111;
        rom_memory[24285] = 3'b111;
        rom_memory[24286] = 3'b111;
        rom_memory[24287] = 3'b111;
        rom_memory[24288] = 3'b111;
        rom_memory[24289] = 3'b111;
        rom_memory[24290] = 3'b111;
        rom_memory[24291] = 3'b111;
        rom_memory[24292] = 3'b110;
        rom_memory[24293] = 3'b100;
        rom_memory[24294] = 3'b110;
        rom_memory[24295] = 3'b110;
        rom_memory[24296] = 3'b100;
        rom_memory[24297] = 3'b100;
        rom_memory[24298] = 3'b100;
        rom_memory[24299] = 3'b100;
        rom_memory[24300] = 3'b100;
        rom_memory[24301] = 3'b100;
        rom_memory[24302] = 3'b100;
        rom_memory[24303] = 3'b110;
        rom_memory[24304] = 3'b110;
        rom_memory[24305] = 3'b110;
        rom_memory[24306] = 3'b110;
        rom_memory[24307] = 3'b110;
        rom_memory[24308] = 3'b110;
        rom_memory[24309] = 3'b110;
        rom_memory[24310] = 3'b110;
        rom_memory[24311] = 3'b110;
        rom_memory[24312] = 3'b110;
        rom_memory[24313] = 3'b110;
        rom_memory[24314] = 3'b110;
        rom_memory[24315] = 3'b110;
        rom_memory[24316] = 3'b110;
        rom_memory[24317] = 3'b110;
        rom_memory[24318] = 3'b110;
        rom_memory[24319] = 3'b110;
        rom_memory[24320] = 3'b110;
        rom_memory[24321] = 3'b110;
        rom_memory[24322] = 3'b110;
        rom_memory[24323] = 3'b110;
        rom_memory[24324] = 3'b110;
        rom_memory[24325] = 3'b110;
        rom_memory[24326] = 3'b110;
        rom_memory[24327] = 3'b110;
        rom_memory[24328] = 3'b110;
        rom_memory[24329] = 3'b110;
        rom_memory[24330] = 3'b110;
        rom_memory[24331] = 3'b110;
        rom_memory[24332] = 3'b110;
        rom_memory[24333] = 3'b110;
        rom_memory[24334] = 3'b110;
        rom_memory[24335] = 3'b110;
        rom_memory[24336] = 3'b110;
        rom_memory[24337] = 3'b110;
        rom_memory[24338] = 3'b110;
        rom_memory[24339] = 3'b110;
        rom_memory[24340] = 3'b110;
        rom_memory[24341] = 3'b110;
        rom_memory[24342] = 3'b110;
        rom_memory[24343] = 3'b110;
        rom_memory[24344] = 3'b110;
        rom_memory[24345] = 3'b110;
        rom_memory[24346] = 3'b111;
        rom_memory[24347] = 3'b111;
        rom_memory[24348] = 3'b111;
        rom_memory[24349] = 3'b111;
        rom_memory[24350] = 3'b111;
        rom_memory[24351] = 3'b111;
        rom_memory[24352] = 3'b111;
        rom_memory[24353] = 3'b111;
        rom_memory[24354] = 3'b111;
        rom_memory[24355] = 3'b111;
        rom_memory[24356] = 3'b111;
        rom_memory[24357] = 3'b110;
        rom_memory[24358] = 3'b000;
        rom_memory[24359] = 3'b000;
        rom_memory[24360] = 3'b000;
        rom_memory[24361] = 3'b000;
        rom_memory[24362] = 3'b000;
        rom_memory[24363] = 3'b000;
        rom_memory[24364] = 3'b000;
        rom_memory[24365] = 3'b000;
        rom_memory[24366] = 3'b000;
        rom_memory[24367] = 3'b000;
        rom_memory[24368] = 3'b110;
        rom_memory[24369] = 3'b110;
        rom_memory[24370] = 3'b110;
        rom_memory[24371] = 3'b110;
        rom_memory[24372] = 3'b110;
        rom_memory[24373] = 3'b110;
        rom_memory[24374] = 3'b110;
        rom_memory[24375] = 3'b110;
        rom_memory[24376] = 3'b110;
        rom_memory[24377] = 3'b110;
        rom_memory[24378] = 3'b110;
        rom_memory[24379] = 3'b110;
        rom_memory[24380] = 3'b110;
        rom_memory[24381] = 3'b110;
        rom_memory[24382] = 3'b110;
        rom_memory[24383] = 3'b110;
        rom_memory[24384] = 3'b110;
        rom_memory[24385] = 3'b110;
        rom_memory[24386] = 3'b110;
        rom_memory[24387] = 3'b110;
        rom_memory[24388] = 3'b110;
        rom_memory[24389] = 3'b110;
        rom_memory[24390] = 3'b110;
        rom_memory[24391] = 3'b110;
        rom_memory[24392] = 3'b110;
        rom_memory[24393] = 3'b110;
        rom_memory[24394] = 3'b110;
        rom_memory[24395] = 3'b110;
        rom_memory[24396] = 3'b110;
        rom_memory[24397] = 3'b110;
        rom_memory[24398] = 3'b110;
        rom_memory[24399] = 3'b110;
        rom_memory[24400] = 3'b110;
        rom_memory[24401] = 3'b110;
        rom_memory[24402] = 3'b110;
        rom_memory[24403] = 3'b110;
        rom_memory[24404] = 3'b111;
        rom_memory[24405] = 3'b111;
        rom_memory[24406] = 3'b111;
        rom_memory[24407] = 3'b111;
        rom_memory[24408] = 3'b111;
        rom_memory[24409] = 3'b111;
        rom_memory[24410] = 3'b110;
        rom_memory[24411] = 3'b111;
        rom_memory[24412] = 3'b111;
        rom_memory[24413] = 3'b111;
        rom_memory[24414] = 3'b111;
        rom_memory[24415] = 3'b111;
        rom_memory[24416] = 3'b111;
        rom_memory[24417] = 3'b111;
        rom_memory[24418] = 3'b111;
        rom_memory[24419] = 3'b111;
        rom_memory[24420] = 3'b111;
        rom_memory[24421] = 3'b111;
        rom_memory[24422] = 3'b111;
        rom_memory[24423] = 3'b111;
        rom_memory[24424] = 3'b110;
        rom_memory[24425] = 3'b110;
        rom_memory[24426] = 3'b111;
        rom_memory[24427] = 3'b111;
        rom_memory[24428] = 3'b111;
        rom_memory[24429] = 3'b111;
        rom_memory[24430] = 3'b111;
        rom_memory[24431] = 3'b111;
        rom_memory[24432] = 3'b111;
        rom_memory[24433] = 3'b111;
        rom_memory[24434] = 3'b111;
        rom_memory[24435] = 3'b111;
        rom_memory[24436] = 3'b111;
        rom_memory[24437] = 3'b111;
        rom_memory[24438] = 3'b111;
        rom_memory[24439] = 3'b111;
        rom_memory[24440] = 3'b111;
        rom_memory[24441] = 3'b111;
        rom_memory[24442] = 3'b111;
        rom_memory[24443] = 3'b111;
        rom_memory[24444] = 3'b111;
        rom_memory[24445] = 3'b111;
        rom_memory[24446] = 3'b111;
        rom_memory[24447] = 3'b111;
        rom_memory[24448] = 3'b111;
        rom_memory[24449] = 3'b111;
        rom_memory[24450] = 3'b111;
        rom_memory[24451] = 3'b111;
        rom_memory[24452] = 3'b111;
        rom_memory[24453] = 3'b111;
        rom_memory[24454] = 3'b111;
        rom_memory[24455] = 3'b111;
        rom_memory[24456] = 3'b111;
        rom_memory[24457] = 3'b111;
        rom_memory[24458] = 3'b111;
        rom_memory[24459] = 3'b111;
        rom_memory[24460] = 3'b111;
        rom_memory[24461] = 3'b111;
        rom_memory[24462] = 3'b111;
        rom_memory[24463] = 3'b111;
        rom_memory[24464] = 3'b111;
        rom_memory[24465] = 3'b111;
        rom_memory[24466] = 3'b111;
        rom_memory[24467] = 3'b111;
        rom_memory[24468] = 3'b111;
        rom_memory[24469] = 3'b111;
        rom_memory[24470] = 3'b111;
        rom_memory[24471] = 3'b111;
        rom_memory[24472] = 3'b111;
        rom_memory[24473] = 3'b111;
        rom_memory[24474] = 3'b111;
        rom_memory[24475] = 3'b111;
        rom_memory[24476] = 3'b111;
        rom_memory[24477] = 3'b111;
        rom_memory[24478] = 3'b111;
        rom_memory[24479] = 3'b111;
        rom_memory[24480] = 3'b110;
        rom_memory[24481] = 3'b110;
        rom_memory[24482] = 3'b110;
        rom_memory[24483] = 3'b110;
        rom_memory[24484] = 3'b110;
        rom_memory[24485] = 3'b110;
        rom_memory[24486] = 3'b110;
        rom_memory[24487] = 3'b110;
        rom_memory[24488] = 3'b110;
        rom_memory[24489] = 3'b110;
        rom_memory[24490] = 3'b110;
        rom_memory[24491] = 3'b110;
        rom_memory[24492] = 3'b110;
        rom_memory[24493] = 3'b110;
        rom_memory[24494] = 3'b110;
        rom_memory[24495] = 3'b110;
        rom_memory[24496] = 3'b110;
        rom_memory[24497] = 3'b110;
        rom_memory[24498] = 3'b110;
        rom_memory[24499] = 3'b110;
        rom_memory[24500] = 3'b110;
        rom_memory[24501] = 3'b110;
        rom_memory[24502] = 3'b110;
        rom_memory[24503] = 3'b110;
        rom_memory[24504] = 3'b110;
        rom_memory[24505] = 3'b110;
        rom_memory[24506] = 3'b110;
        rom_memory[24507] = 3'b110;
        rom_memory[24508] = 3'b111;
        rom_memory[24509] = 3'b111;
        rom_memory[24510] = 3'b111;
        rom_memory[24511] = 3'b111;
        rom_memory[24512] = 3'b111;
        rom_memory[24513] = 3'b111;
        rom_memory[24514] = 3'b111;
        rom_memory[24515] = 3'b111;
        rom_memory[24516] = 3'b111;
        rom_memory[24517] = 3'b111;
        rom_memory[24518] = 3'b111;
        rom_memory[24519] = 3'b111;
        rom_memory[24520] = 3'b111;
        rom_memory[24521] = 3'b111;
        rom_memory[24522] = 3'b111;
        rom_memory[24523] = 3'b111;
        rom_memory[24524] = 3'b111;
        rom_memory[24525] = 3'b111;
        rom_memory[24526] = 3'b111;
        rom_memory[24527] = 3'b111;
        rom_memory[24528] = 3'b111;
        rom_memory[24529] = 3'b111;
        rom_memory[24530] = 3'b111;
        rom_memory[24531] = 3'b111;
        rom_memory[24532] = 3'b110;
        rom_memory[24533] = 3'b110;
        rom_memory[24534] = 3'b100;
        rom_memory[24535] = 3'b110;
        rom_memory[24536] = 3'b100;
        rom_memory[24537] = 3'b100;
        rom_memory[24538] = 3'b100;
        rom_memory[24539] = 3'b100;
        rom_memory[24540] = 3'b100;
        rom_memory[24541] = 3'b100;
        rom_memory[24542] = 3'b100;
        rom_memory[24543] = 3'b110;
        rom_memory[24544] = 3'b110;
        rom_memory[24545] = 3'b110;
        rom_memory[24546] = 3'b110;
        rom_memory[24547] = 3'b110;
        rom_memory[24548] = 3'b110;
        rom_memory[24549] = 3'b110;
        rom_memory[24550] = 3'b110;
        rom_memory[24551] = 3'b110;
        rom_memory[24552] = 3'b110;
        rom_memory[24553] = 3'b110;
        rom_memory[24554] = 3'b110;
        rom_memory[24555] = 3'b110;
        rom_memory[24556] = 3'b110;
        rom_memory[24557] = 3'b110;
        rom_memory[24558] = 3'b110;
        rom_memory[24559] = 3'b110;
        rom_memory[24560] = 3'b110;
        rom_memory[24561] = 3'b110;
        rom_memory[24562] = 3'b110;
        rom_memory[24563] = 3'b110;
        rom_memory[24564] = 3'b110;
        rom_memory[24565] = 3'b110;
        rom_memory[24566] = 3'b110;
        rom_memory[24567] = 3'b110;
        rom_memory[24568] = 3'b110;
        rom_memory[24569] = 3'b110;
        rom_memory[24570] = 3'b110;
        rom_memory[24571] = 3'b110;
        rom_memory[24572] = 3'b110;
        rom_memory[24573] = 3'b110;
        rom_memory[24574] = 3'b110;
        rom_memory[24575] = 3'b110;
        rom_memory[24576] = 3'b110;
        rom_memory[24577] = 3'b110;
        rom_memory[24578] = 3'b110;
        rom_memory[24579] = 3'b110;
        rom_memory[24580] = 3'b110;
        rom_memory[24581] = 3'b110;
        rom_memory[24582] = 3'b110;
        rom_memory[24583] = 3'b110;
        rom_memory[24584] = 3'b110;
        rom_memory[24585] = 3'b110;
        rom_memory[24586] = 3'b111;
        rom_memory[24587] = 3'b110;
        rom_memory[24588] = 3'b110;
        rom_memory[24589] = 3'b111;
        rom_memory[24590] = 3'b111;
        rom_memory[24591] = 3'b111;
        rom_memory[24592] = 3'b111;
        rom_memory[24593] = 3'b111;
        rom_memory[24594] = 3'b111;
        rom_memory[24595] = 3'b111;
        rom_memory[24596] = 3'b111;
        rom_memory[24597] = 3'b110;
        rom_memory[24598] = 3'b100;
        rom_memory[24599] = 3'b000;
        rom_memory[24600] = 3'b000;
        rom_memory[24601] = 3'b000;
        rom_memory[24602] = 3'b000;
        rom_memory[24603] = 3'b000;
        rom_memory[24604] = 3'b000;
        rom_memory[24605] = 3'b000;
        rom_memory[24606] = 3'b000;
        rom_memory[24607] = 3'b000;
        rom_memory[24608] = 3'b000;
        rom_memory[24609] = 3'b110;
        rom_memory[24610] = 3'b110;
        rom_memory[24611] = 3'b110;
        rom_memory[24612] = 3'b110;
        rom_memory[24613] = 3'b110;
        rom_memory[24614] = 3'b110;
        rom_memory[24615] = 3'b110;
        rom_memory[24616] = 3'b110;
        rom_memory[24617] = 3'b110;
        rom_memory[24618] = 3'b110;
        rom_memory[24619] = 3'b110;
        rom_memory[24620] = 3'b110;
        rom_memory[24621] = 3'b110;
        rom_memory[24622] = 3'b110;
        rom_memory[24623] = 3'b110;
        rom_memory[24624] = 3'b110;
        rom_memory[24625] = 3'b110;
        rom_memory[24626] = 3'b110;
        rom_memory[24627] = 3'b110;
        rom_memory[24628] = 3'b110;
        rom_memory[24629] = 3'b110;
        rom_memory[24630] = 3'b110;
        rom_memory[24631] = 3'b110;
        rom_memory[24632] = 3'b110;
        rom_memory[24633] = 3'b110;
        rom_memory[24634] = 3'b110;
        rom_memory[24635] = 3'b110;
        rom_memory[24636] = 3'b110;
        rom_memory[24637] = 3'b110;
        rom_memory[24638] = 3'b110;
        rom_memory[24639] = 3'b110;
        rom_memory[24640] = 3'b110;
        rom_memory[24641] = 3'b110;
        rom_memory[24642] = 3'b110;
        rom_memory[24643] = 3'b110;
        rom_memory[24644] = 3'b110;
        rom_memory[24645] = 3'b110;
        rom_memory[24646] = 3'b110;
        rom_memory[24647] = 3'b110;
        rom_memory[24648] = 3'b111;
        rom_memory[24649] = 3'b111;
        rom_memory[24650] = 3'b111;
        rom_memory[24651] = 3'b111;
        rom_memory[24652] = 3'b111;
        rom_memory[24653] = 3'b111;
        rom_memory[24654] = 3'b111;
        rom_memory[24655] = 3'b111;
        rom_memory[24656] = 3'b111;
        rom_memory[24657] = 3'b111;
        rom_memory[24658] = 3'b111;
        rom_memory[24659] = 3'b111;
        rom_memory[24660] = 3'b111;
        rom_memory[24661] = 3'b111;
        rom_memory[24662] = 3'b111;
        rom_memory[24663] = 3'b111;
        rom_memory[24664] = 3'b111;
        rom_memory[24665] = 3'b111;
        rom_memory[24666] = 3'b111;
        rom_memory[24667] = 3'b111;
        rom_memory[24668] = 3'b111;
        rom_memory[24669] = 3'b111;
        rom_memory[24670] = 3'b111;
        rom_memory[24671] = 3'b111;
        rom_memory[24672] = 3'b111;
        rom_memory[24673] = 3'b111;
        rom_memory[24674] = 3'b111;
        rom_memory[24675] = 3'b111;
        rom_memory[24676] = 3'b111;
        rom_memory[24677] = 3'b111;
        rom_memory[24678] = 3'b111;
        rom_memory[24679] = 3'b111;
        rom_memory[24680] = 3'b111;
        rom_memory[24681] = 3'b111;
        rom_memory[24682] = 3'b111;
        rom_memory[24683] = 3'b111;
        rom_memory[24684] = 3'b111;
        rom_memory[24685] = 3'b111;
        rom_memory[24686] = 3'b111;
        rom_memory[24687] = 3'b111;
        rom_memory[24688] = 3'b111;
        rom_memory[24689] = 3'b111;
        rom_memory[24690] = 3'b111;
        rom_memory[24691] = 3'b111;
        rom_memory[24692] = 3'b111;
        rom_memory[24693] = 3'b111;
        rom_memory[24694] = 3'b111;
        rom_memory[24695] = 3'b111;
        rom_memory[24696] = 3'b111;
        rom_memory[24697] = 3'b111;
        rom_memory[24698] = 3'b111;
        rom_memory[24699] = 3'b111;
        rom_memory[24700] = 3'b111;
        rom_memory[24701] = 3'b111;
        rom_memory[24702] = 3'b111;
        rom_memory[24703] = 3'b111;
        rom_memory[24704] = 3'b111;
        rom_memory[24705] = 3'b111;
        rom_memory[24706] = 3'b111;
        rom_memory[24707] = 3'b111;
        rom_memory[24708] = 3'b111;
        rom_memory[24709] = 3'b111;
        rom_memory[24710] = 3'b111;
        rom_memory[24711] = 3'b111;
        rom_memory[24712] = 3'b111;
        rom_memory[24713] = 3'b111;
        rom_memory[24714] = 3'b111;
        rom_memory[24715] = 3'b111;
        rom_memory[24716] = 3'b111;
        rom_memory[24717] = 3'b111;
        rom_memory[24718] = 3'b111;
        rom_memory[24719] = 3'b111;
        rom_memory[24720] = 3'b110;
        rom_memory[24721] = 3'b110;
        rom_memory[24722] = 3'b110;
        rom_memory[24723] = 3'b110;
        rom_memory[24724] = 3'b110;
        rom_memory[24725] = 3'b110;
        rom_memory[24726] = 3'b110;
        rom_memory[24727] = 3'b110;
        rom_memory[24728] = 3'b110;
        rom_memory[24729] = 3'b110;
        rom_memory[24730] = 3'b110;
        rom_memory[24731] = 3'b110;
        rom_memory[24732] = 3'b110;
        rom_memory[24733] = 3'b110;
        rom_memory[24734] = 3'b110;
        rom_memory[24735] = 3'b110;
        rom_memory[24736] = 3'b110;
        rom_memory[24737] = 3'b110;
        rom_memory[24738] = 3'b110;
        rom_memory[24739] = 3'b110;
        rom_memory[24740] = 3'b110;
        rom_memory[24741] = 3'b110;
        rom_memory[24742] = 3'b110;
        rom_memory[24743] = 3'b110;
        rom_memory[24744] = 3'b110;
        rom_memory[24745] = 3'b110;
        rom_memory[24746] = 3'b110;
        rom_memory[24747] = 3'b110;
        rom_memory[24748] = 3'b111;
        rom_memory[24749] = 3'b111;
        rom_memory[24750] = 3'b111;
        rom_memory[24751] = 3'b111;
        rom_memory[24752] = 3'b111;
        rom_memory[24753] = 3'b111;
        rom_memory[24754] = 3'b111;
        rom_memory[24755] = 3'b111;
        rom_memory[24756] = 3'b111;
        rom_memory[24757] = 3'b111;
        rom_memory[24758] = 3'b111;
        rom_memory[24759] = 3'b111;
        rom_memory[24760] = 3'b111;
        rom_memory[24761] = 3'b111;
        rom_memory[24762] = 3'b111;
        rom_memory[24763] = 3'b111;
        rom_memory[24764] = 3'b111;
        rom_memory[24765] = 3'b111;
        rom_memory[24766] = 3'b111;
        rom_memory[24767] = 3'b111;
        rom_memory[24768] = 3'b111;
        rom_memory[24769] = 3'b111;
        rom_memory[24770] = 3'b111;
        rom_memory[24771] = 3'b111;
        rom_memory[24772] = 3'b111;
        rom_memory[24773] = 3'b110;
        rom_memory[24774] = 3'b100;
        rom_memory[24775] = 3'b110;
        rom_memory[24776] = 3'b100;
        rom_memory[24777] = 3'b100;
        rom_memory[24778] = 3'b100;
        rom_memory[24779] = 3'b100;
        rom_memory[24780] = 3'b100;
        rom_memory[24781] = 3'b100;
        rom_memory[24782] = 3'b100;
        rom_memory[24783] = 3'b100;
        rom_memory[24784] = 3'b100;
        rom_memory[24785] = 3'b110;
        rom_memory[24786] = 3'b110;
        rom_memory[24787] = 3'b110;
        rom_memory[24788] = 3'b110;
        rom_memory[24789] = 3'b110;
        rom_memory[24790] = 3'b110;
        rom_memory[24791] = 3'b110;
        rom_memory[24792] = 3'b110;
        rom_memory[24793] = 3'b110;
        rom_memory[24794] = 3'b110;
        rom_memory[24795] = 3'b110;
        rom_memory[24796] = 3'b110;
        rom_memory[24797] = 3'b110;
        rom_memory[24798] = 3'b110;
        rom_memory[24799] = 3'b110;
        rom_memory[24800] = 3'b110;
        rom_memory[24801] = 3'b110;
        rom_memory[24802] = 3'b110;
        rom_memory[24803] = 3'b110;
        rom_memory[24804] = 3'b110;
        rom_memory[24805] = 3'b110;
        rom_memory[24806] = 3'b110;
        rom_memory[24807] = 3'b110;
        rom_memory[24808] = 3'b110;
        rom_memory[24809] = 3'b110;
        rom_memory[24810] = 3'b110;
        rom_memory[24811] = 3'b110;
        rom_memory[24812] = 3'b110;
        rom_memory[24813] = 3'b110;
        rom_memory[24814] = 3'b110;
        rom_memory[24815] = 3'b110;
        rom_memory[24816] = 3'b110;
        rom_memory[24817] = 3'b110;
        rom_memory[24818] = 3'b110;
        rom_memory[24819] = 3'b110;
        rom_memory[24820] = 3'b110;
        rom_memory[24821] = 3'b110;
        rom_memory[24822] = 3'b110;
        rom_memory[24823] = 3'b110;
        rom_memory[24824] = 3'b110;
        rom_memory[24825] = 3'b110;
        rom_memory[24826] = 3'b110;
        rom_memory[24827] = 3'b111;
        rom_memory[24828] = 3'b110;
        rom_memory[24829] = 3'b110;
        rom_memory[24830] = 3'b111;
        rom_memory[24831] = 3'b111;
        rom_memory[24832] = 3'b111;
        rom_memory[24833] = 3'b111;
        rom_memory[24834] = 3'b111;
        rom_memory[24835] = 3'b111;
        rom_memory[24836] = 3'b111;
        rom_memory[24837] = 3'b110;
        rom_memory[24838] = 3'b110;
        rom_memory[24839] = 3'b000;
        rom_memory[24840] = 3'b000;
        rom_memory[24841] = 3'b000;
        rom_memory[24842] = 3'b000;
        rom_memory[24843] = 3'b000;
        rom_memory[24844] = 3'b000;
        rom_memory[24845] = 3'b000;
        rom_memory[24846] = 3'b000;
        rom_memory[24847] = 3'b000;
        rom_memory[24848] = 3'b000;
        rom_memory[24849] = 3'b110;
        rom_memory[24850] = 3'b110;
        rom_memory[24851] = 3'b110;
        rom_memory[24852] = 3'b110;
        rom_memory[24853] = 3'b110;
        rom_memory[24854] = 3'b110;
        rom_memory[24855] = 3'b110;
        rom_memory[24856] = 3'b110;
        rom_memory[24857] = 3'b110;
        rom_memory[24858] = 3'b110;
        rom_memory[24859] = 3'b110;
        rom_memory[24860] = 3'b110;
        rom_memory[24861] = 3'b110;
        rom_memory[24862] = 3'b110;
        rom_memory[24863] = 3'b110;
        rom_memory[24864] = 3'b110;
        rom_memory[24865] = 3'b110;
        rom_memory[24866] = 3'b110;
        rom_memory[24867] = 3'b110;
        rom_memory[24868] = 3'b110;
        rom_memory[24869] = 3'b110;
        rom_memory[24870] = 3'b110;
        rom_memory[24871] = 3'b110;
        rom_memory[24872] = 3'b110;
        rom_memory[24873] = 3'b110;
        rom_memory[24874] = 3'b110;
        rom_memory[24875] = 3'b110;
        rom_memory[24876] = 3'b110;
        rom_memory[24877] = 3'b110;
        rom_memory[24878] = 3'b110;
        rom_memory[24879] = 3'b110;
        rom_memory[24880] = 3'b110;
        rom_memory[24881] = 3'b110;
        rom_memory[24882] = 3'b110;
        rom_memory[24883] = 3'b110;
        rom_memory[24884] = 3'b110;
        rom_memory[24885] = 3'b111;
        rom_memory[24886] = 3'b111;
        rom_memory[24887] = 3'b110;
        rom_memory[24888] = 3'b110;
        rom_memory[24889] = 3'b111;
        rom_memory[24890] = 3'b111;
        rom_memory[24891] = 3'b111;
        rom_memory[24892] = 3'b111;
        rom_memory[24893] = 3'b111;
        rom_memory[24894] = 3'b111;
        rom_memory[24895] = 3'b111;
        rom_memory[24896] = 3'b111;
        rom_memory[24897] = 3'b111;
        rom_memory[24898] = 3'b111;
        rom_memory[24899] = 3'b111;
        rom_memory[24900] = 3'b111;
        rom_memory[24901] = 3'b111;
        rom_memory[24902] = 3'b111;
        rom_memory[24903] = 3'b111;
        rom_memory[24904] = 3'b111;
        rom_memory[24905] = 3'b111;
        rom_memory[24906] = 3'b111;
        rom_memory[24907] = 3'b111;
        rom_memory[24908] = 3'b111;
        rom_memory[24909] = 3'b111;
        rom_memory[24910] = 3'b111;
        rom_memory[24911] = 3'b111;
        rom_memory[24912] = 3'b111;
        rom_memory[24913] = 3'b111;
        rom_memory[24914] = 3'b111;
        rom_memory[24915] = 3'b111;
        rom_memory[24916] = 3'b111;
        rom_memory[24917] = 3'b111;
        rom_memory[24918] = 3'b111;
        rom_memory[24919] = 3'b111;
        rom_memory[24920] = 3'b111;
        rom_memory[24921] = 3'b111;
        rom_memory[24922] = 3'b111;
        rom_memory[24923] = 3'b111;
        rom_memory[24924] = 3'b111;
        rom_memory[24925] = 3'b111;
        rom_memory[24926] = 3'b111;
        rom_memory[24927] = 3'b111;
        rom_memory[24928] = 3'b111;
        rom_memory[24929] = 3'b111;
        rom_memory[24930] = 3'b111;
        rom_memory[24931] = 3'b111;
        rom_memory[24932] = 3'b111;
        rom_memory[24933] = 3'b111;
        rom_memory[24934] = 3'b111;
        rom_memory[24935] = 3'b111;
        rom_memory[24936] = 3'b111;
        rom_memory[24937] = 3'b111;
        rom_memory[24938] = 3'b111;
        rom_memory[24939] = 3'b111;
        rom_memory[24940] = 3'b111;
        rom_memory[24941] = 3'b111;
        rom_memory[24942] = 3'b111;
        rom_memory[24943] = 3'b111;
        rom_memory[24944] = 3'b111;
        rom_memory[24945] = 3'b111;
        rom_memory[24946] = 3'b111;
        rom_memory[24947] = 3'b111;
        rom_memory[24948] = 3'b111;
        rom_memory[24949] = 3'b111;
        rom_memory[24950] = 3'b111;
        rom_memory[24951] = 3'b111;
        rom_memory[24952] = 3'b111;
        rom_memory[24953] = 3'b111;
        rom_memory[24954] = 3'b111;
        rom_memory[24955] = 3'b111;
        rom_memory[24956] = 3'b111;
        rom_memory[24957] = 3'b111;
        rom_memory[24958] = 3'b111;
        rom_memory[24959] = 3'b111;
        rom_memory[24960] = 3'b110;
        rom_memory[24961] = 3'b110;
        rom_memory[24962] = 3'b110;
        rom_memory[24963] = 3'b110;
        rom_memory[24964] = 3'b110;
        rom_memory[24965] = 3'b110;
        rom_memory[24966] = 3'b110;
        rom_memory[24967] = 3'b110;
        rom_memory[24968] = 3'b110;
        rom_memory[24969] = 3'b110;
        rom_memory[24970] = 3'b110;
        rom_memory[24971] = 3'b110;
        rom_memory[24972] = 3'b110;
        rom_memory[24973] = 3'b110;
        rom_memory[24974] = 3'b110;
        rom_memory[24975] = 3'b110;
        rom_memory[24976] = 3'b110;
        rom_memory[24977] = 3'b110;
        rom_memory[24978] = 3'b110;
        rom_memory[24979] = 3'b110;
        rom_memory[24980] = 3'b110;
        rom_memory[24981] = 3'b110;
        rom_memory[24982] = 3'b110;
        rom_memory[24983] = 3'b110;
        rom_memory[24984] = 3'b110;
        rom_memory[24985] = 3'b110;
        rom_memory[24986] = 3'b110;
        rom_memory[24987] = 3'b110;
        rom_memory[24988] = 3'b111;
        rom_memory[24989] = 3'b111;
        rom_memory[24990] = 3'b111;
        rom_memory[24991] = 3'b111;
        rom_memory[24992] = 3'b111;
        rom_memory[24993] = 3'b111;
        rom_memory[24994] = 3'b111;
        rom_memory[24995] = 3'b111;
        rom_memory[24996] = 3'b111;
        rom_memory[24997] = 3'b111;
        rom_memory[24998] = 3'b111;
        rom_memory[24999] = 3'b111;
        rom_memory[25000] = 3'b111;
        rom_memory[25001] = 3'b111;
        rom_memory[25002] = 3'b111;
        rom_memory[25003] = 3'b111;
        rom_memory[25004] = 3'b111;
        rom_memory[25005] = 3'b111;
        rom_memory[25006] = 3'b111;
        rom_memory[25007] = 3'b111;
        rom_memory[25008] = 3'b111;
        rom_memory[25009] = 3'b111;
        rom_memory[25010] = 3'b111;
        rom_memory[25011] = 3'b111;
        rom_memory[25012] = 3'b111;
        rom_memory[25013] = 3'b110;
        rom_memory[25014] = 3'b110;
        rom_memory[25015] = 3'b110;
        rom_memory[25016] = 3'b110;
        rom_memory[25017] = 3'b100;
        rom_memory[25018] = 3'b100;
        rom_memory[25019] = 3'b100;
        rom_memory[25020] = 3'b100;
        rom_memory[25021] = 3'b100;
        rom_memory[25022] = 3'b100;
        rom_memory[25023] = 3'b100;
        rom_memory[25024] = 3'b100;
        rom_memory[25025] = 3'b110;
        rom_memory[25026] = 3'b110;
        rom_memory[25027] = 3'b110;
        rom_memory[25028] = 3'b110;
        rom_memory[25029] = 3'b110;
        rom_memory[25030] = 3'b110;
        rom_memory[25031] = 3'b110;
        rom_memory[25032] = 3'b110;
        rom_memory[25033] = 3'b110;
        rom_memory[25034] = 3'b110;
        rom_memory[25035] = 3'b110;
        rom_memory[25036] = 3'b110;
        rom_memory[25037] = 3'b110;
        rom_memory[25038] = 3'b110;
        rom_memory[25039] = 3'b110;
        rom_memory[25040] = 3'b110;
        rom_memory[25041] = 3'b110;
        rom_memory[25042] = 3'b110;
        rom_memory[25043] = 3'b110;
        rom_memory[25044] = 3'b110;
        rom_memory[25045] = 3'b110;
        rom_memory[25046] = 3'b110;
        rom_memory[25047] = 3'b110;
        rom_memory[25048] = 3'b110;
        rom_memory[25049] = 3'b110;
        rom_memory[25050] = 3'b110;
        rom_memory[25051] = 3'b110;
        rom_memory[25052] = 3'b110;
        rom_memory[25053] = 3'b110;
        rom_memory[25054] = 3'b110;
        rom_memory[25055] = 3'b110;
        rom_memory[25056] = 3'b110;
        rom_memory[25057] = 3'b110;
        rom_memory[25058] = 3'b110;
        rom_memory[25059] = 3'b110;
        rom_memory[25060] = 3'b110;
        rom_memory[25061] = 3'b110;
        rom_memory[25062] = 3'b110;
        rom_memory[25063] = 3'b110;
        rom_memory[25064] = 3'b110;
        rom_memory[25065] = 3'b110;
        rom_memory[25066] = 3'b110;
        rom_memory[25067] = 3'b110;
        rom_memory[25068] = 3'b110;
        rom_memory[25069] = 3'b110;
        rom_memory[25070] = 3'b111;
        rom_memory[25071] = 3'b111;
        rom_memory[25072] = 3'b111;
        rom_memory[25073] = 3'b111;
        rom_memory[25074] = 3'b111;
        rom_memory[25075] = 3'b111;
        rom_memory[25076] = 3'b111;
        rom_memory[25077] = 3'b111;
        rom_memory[25078] = 3'b110;
        rom_memory[25079] = 3'b100;
        rom_memory[25080] = 3'b000;
        rom_memory[25081] = 3'b000;
        rom_memory[25082] = 3'b000;
        rom_memory[25083] = 3'b000;
        rom_memory[25084] = 3'b000;
        rom_memory[25085] = 3'b000;
        rom_memory[25086] = 3'b000;
        rom_memory[25087] = 3'b000;
        rom_memory[25088] = 3'b000;
        rom_memory[25089] = 3'b000;
        rom_memory[25090] = 3'b110;
        rom_memory[25091] = 3'b110;
        rom_memory[25092] = 3'b110;
        rom_memory[25093] = 3'b110;
        rom_memory[25094] = 3'b110;
        rom_memory[25095] = 3'b110;
        rom_memory[25096] = 3'b110;
        rom_memory[25097] = 3'b110;
        rom_memory[25098] = 3'b110;
        rom_memory[25099] = 3'b110;
        rom_memory[25100] = 3'b110;
        rom_memory[25101] = 3'b110;
        rom_memory[25102] = 3'b110;
        rom_memory[25103] = 3'b110;
        rom_memory[25104] = 3'b110;
        rom_memory[25105] = 3'b110;
        rom_memory[25106] = 3'b110;
        rom_memory[25107] = 3'b110;
        rom_memory[25108] = 3'b110;
        rom_memory[25109] = 3'b110;
        rom_memory[25110] = 3'b110;
        rom_memory[25111] = 3'b110;
        rom_memory[25112] = 3'b110;
        rom_memory[25113] = 3'b110;
        rom_memory[25114] = 3'b110;
        rom_memory[25115] = 3'b110;
        rom_memory[25116] = 3'b110;
        rom_memory[25117] = 3'b110;
        rom_memory[25118] = 3'b110;
        rom_memory[25119] = 3'b110;
        rom_memory[25120] = 3'b110;
        rom_memory[25121] = 3'b110;
        rom_memory[25122] = 3'b110;
        rom_memory[25123] = 3'b110;
        rom_memory[25124] = 3'b110;
        rom_memory[25125] = 3'b110;
        rom_memory[25126] = 3'b110;
        rom_memory[25127] = 3'b110;
        rom_memory[25128] = 3'b110;
        rom_memory[25129] = 3'b110;
        rom_memory[25130] = 3'b111;
        rom_memory[25131] = 3'b111;
        rom_memory[25132] = 3'b111;
        rom_memory[25133] = 3'b111;
        rom_memory[25134] = 3'b111;
        rom_memory[25135] = 3'b111;
        rom_memory[25136] = 3'b111;
        rom_memory[25137] = 3'b111;
        rom_memory[25138] = 3'b111;
        rom_memory[25139] = 3'b111;
        rom_memory[25140] = 3'b111;
        rom_memory[25141] = 3'b111;
        rom_memory[25142] = 3'b111;
        rom_memory[25143] = 3'b111;
        rom_memory[25144] = 3'b111;
        rom_memory[25145] = 3'b111;
        rom_memory[25146] = 3'b111;
        rom_memory[25147] = 3'b111;
        rom_memory[25148] = 3'b111;
        rom_memory[25149] = 3'b111;
        rom_memory[25150] = 3'b111;
        rom_memory[25151] = 3'b111;
        rom_memory[25152] = 3'b111;
        rom_memory[25153] = 3'b111;
        rom_memory[25154] = 3'b111;
        rom_memory[25155] = 3'b111;
        rom_memory[25156] = 3'b111;
        rom_memory[25157] = 3'b111;
        rom_memory[25158] = 3'b111;
        rom_memory[25159] = 3'b111;
        rom_memory[25160] = 3'b111;
        rom_memory[25161] = 3'b111;
        rom_memory[25162] = 3'b111;
        rom_memory[25163] = 3'b111;
        rom_memory[25164] = 3'b111;
        rom_memory[25165] = 3'b111;
        rom_memory[25166] = 3'b111;
        rom_memory[25167] = 3'b111;
        rom_memory[25168] = 3'b111;
        rom_memory[25169] = 3'b111;
        rom_memory[25170] = 3'b111;
        rom_memory[25171] = 3'b111;
        rom_memory[25172] = 3'b111;
        rom_memory[25173] = 3'b111;
        rom_memory[25174] = 3'b111;
        rom_memory[25175] = 3'b111;
        rom_memory[25176] = 3'b111;
        rom_memory[25177] = 3'b111;
        rom_memory[25178] = 3'b111;
        rom_memory[25179] = 3'b111;
        rom_memory[25180] = 3'b111;
        rom_memory[25181] = 3'b111;
        rom_memory[25182] = 3'b111;
        rom_memory[25183] = 3'b111;
        rom_memory[25184] = 3'b111;
        rom_memory[25185] = 3'b111;
        rom_memory[25186] = 3'b111;
        rom_memory[25187] = 3'b111;
        rom_memory[25188] = 3'b111;
        rom_memory[25189] = 3'b111;
        rom_memory[25190] = 3'b111;
        rom_memory[25191] = 3'b111;
        rom_memory[25192] = 3'b111;
        rom_memory[25193] = 3'b111;
        rom_memory[25194] = 3'b111;
        rom_memory[25195] = 3'b111;
        rom_memory[25196] = 3'b111;
        rom_memory[25197] = 3'b111;
        rom_memory[25198] = 3'b111;
        rom_memory[25199] = 3'b111;
        rom_memory[25200] = 3'b110;
        rom_memory[25201] = 3'b110;
        rom_memory[25202] = 3'b110;
        rom_memory[25203] = 3'b110;
        rom_memory[25204] = 3'b110;
        rom_memory[25205] = 3'b110;
        rom_memory[25206] = 3'b110;
        rom_memory[25207] = 3'b110;
        rom_memory[25208] = 3'b110;
        rom_memory[25209] = 3'b110;
        rom_memory[25210] = 3'b110;
        rom_memory[25211] = 3'b110;
        rom_memory[25212] = 3'b110;
        rom_memory[25213] = 3'b110;
        rom_memory[25214] = 3'b110;
        rom_memory[25215] = 3'b110;
        rom_memory[25216] = 3'b110;
        rom_memory[25217] = 3'b110;
        rom_memory[25218] = 3'b110;
        rom_memory[25219] = 3'b110;
        rom_memory[25220] = 3'b110;
        rom_memory[25221] = 3'b110;
        rom_memory[25222] = 3'b110;
        rom_memory[25223] = 3'b110;
        rom_memory[25224] = 3'b110;
        rom_memory[25225] = 3'b110;
        rom_memory[25226] = 3'b110;
        rom_memory[25227] = 3'b110;
        rom_memory[25228] = 3'b111;
        rom_memory[25229] = 3'b111;
        rom_memory[25230] = 3'b111;
        rom_memory[25231] = 3'b111;
        rom_memory[25232] = 3'b111;
        rom_memory[25233] = 3'b111;
        rom_memory[25234] = 3'b111;
        rom_memory[25235] = 3'b111;
        rom_memory[25236] = 3'b111;
        rom_memory[25237] = 3'b111;
        rom_memory[25238] = 3'b111;
        rom_memory[25239] = 3'b111;
        rom_memory[25240] = 3'b111;
        rom_memory[25241] = 3'b111;
        rom_memory[25242] = 3'b111;
        rom_memory[25243] = 3'b111;
        rom_memory[25244] = 3'b111;
        rom_memory[25245] = 3'b111;
        rom_memory[25246] = 3'b111;
        rom_memory[25247] = 3'b111;
        rom_memory[25248] = 3'b111;
        rom_memory[25249] = 3'b111;
        rom_memory[25250] = 3'b111;
        rom_memory[25251] = 3'b111;
        rom_memory[25252] = 3'b111;
        rom_memory[25253] = 3'b111;
        rom_memory[25254] = 3'b110;
        rom_memory[25255] = 3'b110;
        rom_memory[25256] = 3'b110;
        rom_memory[25257] = 3'b100;
        rom_memory[25258] = 3'b110;
        rom_memory[25259] = 3'b110;
        rom_memory[25260] = 3'b100;
        rom_memory[25261] = 3'b100;
        rom_memory[25262] = 3'b100;
        rom_memory[25263] = 3'b100;
        rom_memory[25264] = 3'b100;
        rom_memory[25265] = 3'b100;
        rom_memory[25266] = 3'b110;
        rom_memory[25267] = 3'b110;
        rom_memory[25268] = 3'b110;
        rom_memory[25269] = 3'b110;
        rom_memory[25270] = 3'b110;
        rom_memory[25271] = 3'b110;
        rom_memory[25272] = 3'b110;
        rom_memory[25273] = 3'b110;
        rom_memory[25274] = 3'b110;
        rom_memory[25275] = 3'b110;
        rom_memory[25276] = 3'b110;
        rom_memory[25277] = 3'b110;
        rom_memory[25278] = 3'b110;
        rom_memory[25279] = 3'b110;
        rom_memory[25280] = 3'b110;
        rom_memory[25281] = 3'b110;
        rom_memory[25282] = 3'b110;
        rom_memory[25283] = 3'b110;
        rom_memory[25284] = 3'b110;
        rom_memory[25285] = 3'b110;
        rom_memory[25286] = 3'b110;
        rom_memory[25287] = 3'b110;
        rom_memory[25288] = 3'b110;
        rom_memory[25289] = 3'b110;
        rom_memory[25290] = 3'b110;
        rom_memory[25291] = 3'b110;
        rom_memory[25292] = 3'b110;
        rom_memory[25293] = 3'b110;
        rom_memory[25294] = 3'b110;
        rom_memory[25295] = 3'b110;
        rom_memory[25296] = 3'b110;
        rom_memory[25297] = 3'b110;
        rom_memory[25298] = 3'b110;
        rom_memory[25299] = 3'b110;
        rom_memory[25300] = 3'b110;
        rom_memory[25301] = 3'b110;
        rom_memory[25302] = 3'b110;
        rom_memory[25303] = 3'b110;
        rom_memory[25304] = 3'b110;
        rom_memory[25305] = 3'b110;
        rom_memory[25306] = 3'b110;
        rom_memory[25307] = 3'b110;
        rom_memory[25308] = 3'b110;
        rom_memory[25309] = 3'b110;
        rom_memory[25310] = 3'b110;
        rom_memory[25311] = 3'b111;
        rom_memory[25312] = 3'b111;
        rom_memory[25313] = 3'b110;
        rom_memory[25314] = 3'b110;
        rom_memory[25315] = 3'b111;
        rom_memory[25316] = 3'b111;
        rom_memory[25317] = 3'b111;
        rom_memory[25318] = 3'b110;
        rom_memory[25319] = 3'b110;
        rom_memory[25320] = 3'b000;
        rom_memory[25321] = 3'b000;
        rom_memory[25322] = 3'b000;
        rom_memory[25323] = 3'b000;
        rom_memory[25324] = 3'b000;
        rom_memory[25325] = 3'b000;
        rom_memory[25326] = 3'b000;
        rom_memory[25327] = 3'b000;
        rom_memory[25328] = 3'b000;
        rom_memory[25329] = 3'b000;
        rom_memory[25330] = 3'b000;
        rom_memory[25331] = 3'b110;
        rom_memory[25332] = 3'b110;
        rom_memory[25333] = 3'b110;
        rom_memory[25334] = 3'b110;
        rom_memory[25335] = 3'b110;
        rom_memory[25336] = 3'b110;
        rom_memory[25337] = 3'b110;
        rom_memory[25338] = 3'b110;
        rom_memory[25339] = 3'b110;
        rom_memory[25340] = 3'b110;
        rom_memory[25341] = 3'b110;
        rom_memory[25342] = 3'b110;
        rom_memory[25343] = 3'b110;
        rom_memory[25344] = 3'b110;
        rom_memory[25345] = 3'b110;
        rom_memory[25346] = 3'b110;
        rom_memory[25347] = 3'b110;
        rom_memory[25348] = 3'b110;
        rom_memory[25349] = 3'b110;
        rom_memory[25350] = 3'b110;
        rom_memory[25351] = 3'b110;
        rom_memory[25352] = 3'b110;
        rom_memory[25353] = 3'b110;
        rom_memory[25354] = 3'b110;
        rom_memory[25355] = 3'b110;
        rom_memory[25356] = 3'b110;
        rom_memory[25357] = 3'b110;
        rom_memory[25358] = 3'b110;
        rom_memory[25359] = 3'b110;
        rom_memory[25360] = 3'b110;
        rom_memory[25361] = 3'b110;
        rom_memory[25362] = 3'b110;
        rom_memory[25363] = 3'b110;
        rom_memory[25364] = 3'b110;
        rom_memory[25365] = 3'b110;
        rom_memory[25366] = 3'b111;
        rom_memory[25367] = 3'b110;
        rom_memory[25368] = 3'b110;
        rom_memory[25369] = 3'b110;
        rom_memory[25370] = 3'b111;
        rom_memory[25371] = 3'b111;
        rom_memory[25372] = 3'b111;
        rom_memory[25373] = 3'b111;
        rom_memory[25374] = 3'b111;
        rom_memory[25375] = 3'b111;
        rom_memory[25376] = 3'b111;
        rom_memory[25377] = 3'b111;
        rom_memory[25378] = 3'b111;
        rom_memory[25379] = 3'b111;
        rom_memory[25380] = 3'b111;
        rom_memory[25381] = 3'b111;
        rom_memory[25382] = 3'b111;
        rom_memory[25383] = 3'b111;
        rom_memory[25384] = 3'b111;
        rom_memory[25385] = 3'b111;
        rom_memory[25386] = 3'b111;
        rom_memory[25387] = 3'b111;
        rom_memory[25388] = 3'b111;
        rom_memory[25389] = 3'b111;
        rom_memory[25390] = 3'b111;
        rom_memory[25391] = 3'b111;
        rom_memory[25392] = 3'b111;
        rom_memory[25393] = 3'b111;
        rom_memory[25394] = 3'b111;
        rom_memory[25395] = 3'b111;
        rom_memory[25396] = 3'b111;
        rom_memory[25397] = 3'b111;
        rom_memory[25398] = 3'b111;
        rom_memory[25399] = 3'b111;
        rom_memory[25400] = 3'b111;
        rom_memory[25401] = 3'b111;
        rom_memory[25402] = 3'b111;
        rom_memory[25403] = 3'b111;
        rom_memory[25404] = 3'b111;
        rom_memory[25405] = 3'b111;
        rom_memory[25406] = 3'b111;
        rom_memory[25407] = 3'b111;
        rom_memory[25408] = 3'b111;
        rom_memory[25409] = 3'b111;
        rom_memory[25410] = 3'b111;
        rom_memory[25411] = 3'b111;
        rom_memory[25412] = 3'b111;
        rom_memory[25413] = 3'b111;
        rom_memory[25414] = 3'b111;
        rom_memory[25415] = 3'b111;
        rom_memory[25416] = 3'b111;
        rom_memory[25417] = 3'b111;
        rom_memory[25418] = 3'b111;
        rom_memory[25419] = 3'b111;
        rom_memory[25420] = 3'b111;
        rom_memory[25421] = 3'b111;
        rom_memory[25422] = 3'b111;
        rom_memory[25423] = 3'b111;
        rom_memory[25424] = 3'b111;
        rom_memory[25425] = 3'b111;
        rom_memory[25426] = 3'b111;
        rom_memory[25427] = 3'b111;
        rom_memory[25428] = 3'b111;
        rom_memory[25429] = 3'b111;
        rom_memory[25430] = 3'b111;
        rom_memory[25431] = 3'b111;
        rom_memory[25432] = 3'b111;
        rom_memory[25433] = 3'b111;
        rom_memory[25434] = 3'b111;
        rom_memory[25435] = 3'b111;
        rom_memory[25436] = 3'b111;
        rom_memory[25437] = 3'b111;
        rom_memory[25438] = 3'b111;
        rom_memory[25439] = 3'b111;
        rom_memory[25440] = 3'b110;
        rom_memory[25441] = 3'b110;
        rom_memory[25442] = 3'b110;
        rom_memory[25443] = 3'b110;
        rom_memory[25444] = 3'b110;
        rom_memory[25445] = 3'b110;
        rom_memory[25446] = 3'b110;
        rom_memory[25447] = 3'b110;
        rom_memory[25448] = 3'b110;
        rom_memory[25449] = 3'b110;
        rom_memory[25450] = 3'b110;
        rom_memory[25451] = 3'b110;
        rom_memory[25452] = 3'b110;
        rom_memory[25453] = 3'b110;
        rom_memory[25454] = 3'b110;
        rom_memory[25455] = 3'b110;
        rom_memory[25456] = 3'b110;
        rom_memory[25457] = 3'b110;
        rom_memory[25458] = 3'b110;
        rom_memory[25459] = 3'b110;
        rom_memory[25460] = 3'b110;
        rom_memory[25461] = 3'b110;
        rom_memory[25462] = 3'b110;
        rom_memory[25463] = 3'b110;
        rom_memory[25464] = 3'b110;
        rom_memory[25465] = 3'b110;
        rom_memory[25466] = 3'b110;
        rom_memory[25467] = 3'b110;
        rom_memory[25468] = 3'b110;
        rom_memory[25469] = 3'b111;
        rom_memory[25470] = 3'b111;
        rom_memory[25471] = 3'b111;
        rom_memory[25472] = 3'b111;
        rom_memory[25473] = 3'b111;
        rom_memory[25474] = 3'b111;
        rom_memory[25475] = 3'b111;
        rom_memory[25476] = 3'b111;
        rom_memory[25477] = 3'b111;
        rom_memory[25478] = 3'b111;
        rom_memory[25479] = 3'b111;
        rom_memory[25480] = 3'b111;
        rom_memory[25481] = 3'b111;
        rom_memory[25482] = 3'b111;
        rom_memory[25483] = 3'b111;
        rom_memory[25484] = 3'b111;
        rom_memory[25485] = 3'b111;
        rom_memory[25486] = 3'b111;
        rom_memory[25487] = 3'b111;
        rom_memory[25488] = 3'b111;
        rom_memory[25489] = 3'b111;
        rom_memory[25490] = 3'b111;
        rom_memory[25491] = 3'b111;
        rom_memory[25492] = 3'b111;
        rom_memory[25493] = 3'b111;
        rom_memory[25494] = 3'b111;
        rom_memory[25495] = 3'b110;
        rom_memory[25496] = 3'b110;
        rom_memory[25497] = 3'b110;
        rom_memory[25498] = 3'b110;
        rom_memory[25499] = 3'b110;
        rom_memory[25500] = 3'b110;
        rom_memory[25501] = 3'b100;
        rom_memory[25502] = 3'b100;
        rom_memory[25503] = 3'b100;
        rom_memory[25504] = 3'b100;
        rom_memory[25505] = 3'b100;
        rom_memory[25506] = 3'b100;
        rom_memory[25507] = 3'b100;
        rom_memory[25508] = 3'b110;
        rom_memory[25509] = 3'b110;
        rom_memory[25510] = 3'b110;
        rom_memory[25511] = 3'b110;
        rom_memory[25512] = 3'b110;
        rom_memory[25513] = 3'b110;
        rom_memory[25514] = 3'b110;
        rom_memory[25515] = 3'b110;
        rom_memory[25516] = 3'b110;
        rom_memory[25517] = 3'b110;
        rom_memory[25518] = 3'b110;
        rom_memory[25519] = 3'b110;
        rom_memory[25520] = 3'b110;
        rom_memory[25521] = 3'b110;
        rom_memory[25522] = 3'b110;
        rom_memory[25523] = 3'b110;
        rom_memory[25524] = 3'b110;
        rom_memory[25525] = 3'b110;
        rom_memory[25526] = 3'b110;
        rom_memory[25527] = 3'b110;
        rom_memory[25528] = 3'b110;
        rom_memory[25529] = 3'b110;
        rom_memory[25530] = 3'b110;
        rom_memory[25531] = 3'b110;
        rom_memory[25532] = 3'b110;
        rom_memory[25533] = 3'b110;
        rom_memory[25534] = 3'b110;
        rom_memory[25535] = 3'b110;
        rom_memory[25536] = 3'b110;
        rom_memory[25537] = 3'b110;
        rom_memory[25538] = 3'b110;
        rom_memory[25539] = 3'b110;
        rom_memory[25540] = 3'b110;
        rom_memory[25541] = 3'b110;
        rom_memory[25542] = 3'b110;
        rom_memory[25543] = 3'b110;
        rom_memory[25544] = 3'b110;
        rom_memory[25545] = 3'b110;
        rom_memory[25546] = 3'b110;
        rom_memory[25547] = 3'b110;
        rom_memory[25548] = 3'b110;
        rom_memory[25549] = 3'b110;
        rom_memory[25550] = 3'b110;
        rom_memory[25551] = 3'b110;
        rom_memory[25552] = 3'b111;
        rom_memory[25553] = 3'b110;
        rom_memory[25554] = 3'b110;
        rom_memory[25555] = 3'b110;
        rom_memory[25556] = 3'b110;
        rom_memory[25557] = 3'b110;
        rom_memory[25558] = 3'b110;
        rom_memory[25559] = 3'b110;
        rom_memory[25560] = 3'b000;
        rom_memory[25561] = 3'b000;
        rom_memory[25562] = 3'b000;
        rom_memory[25563] = 3'b000;
        rom_memory[25564] = 3'b000;
        rom_memory[25565] = 3'b000;
        rom_memory[25566] = 3'b000;
        rom_memory[25567] = 3'b000;
        rom_memory[25568] = 3'b000;
        rom_memory[25569] = 3'b000;
        rom_memory[25570] = 3'b000;
        rom_memory[25571] = 3'b110;
        rom_memory[25572] = 3'b110;
        rom_memory[25573] = 3'b110;
        rom_memory[25574] = 3'b110;
        rom_memory[25575] = 3'b110;
        rom_memory[25576] = 3'b110;
        rom_memory[25577] = 3'b110;
        rom_memory[25578] = 3'b110;
        rom_memory[25579] = 3'b110;
        rom_memory[25580] = 3'b110;
        rom_memory[25581] = 3'b110;
        rom_memory[25582] = 3'b110;
        rom_memory[25583] = 3'b110;
        rom_memory[25584] = 3'b110;
        rom_memory[25585] = 3'b110;
        rom_memory[25586] = 3'b110;
        rom_memory[25587] = 3'b110;
        rom_memory[25588] = 3'b110;
        rom_memory[25589] = 3'b110;
        rom_memory[25590] = 3'b110;
        rom_memory[25591] = 3'b110;
        rom_memory[25592] = 3'b110;
        rom_memory[25593] = 3'b110;
        rom_memory[25594] = 3'b110;
        rom_memory[25595] = 3'b110;
        rom_memory[25596] = 3'b110;
        rom_memory[25597] = 3'b110;
        rom_memory[25598] = 3'b110;
        rom_memory[25599] = 3'b110;
        rom_memory[25600] = 3'b110;
        rom_memory[25601] = 3'b110;
        rom_memory[25602] = 3'b110;
        rom_memory[25603] = 3'b110;
        rom_memory[25604] = 3'b110;
        rom_memory[25605] = 3'b110;
        rom_memory[25606] = 3'b110;
        rom_memory[25607] = 3'b110;
        rom_memory[25608] = 3'b110;
        rom_memory[25609] = 3'b110;
        rom_memory[25610] = 3'b111;
        rom_memory[25611] = 3'b111;
        rom_memory[25612] = 3'b111;
        rom_memory[25613] = 3'b111;
        rom_memory[25614] = 3'b111;
        rom_memory[25615] = 3'b111;
        rom_memory[25616] = 3'b111;
        rom_memory[25617] = 3'b111;
        rom_memory[25618] = 3'b111;
        rom_memory[25619] = 3'b111;
        rom_memory[25620] = 3'b111;
        rom_memory[25621] = 3'b111;
        rom_memory[25622] = 3'b111;
        rom_memory[25623] = 3'b111;
        rom_memory[25624] = 3'b111;
        rom_memory[25625] = 3'b111;
        rom_memory[25626] = 3'b111;
        rom_memory[25627] = 3'b111;
        rom_memory[25628] = 3'b111;
        rom_memory[25629] = 3'b111;
        rom_memory[25630] = 3'b111;
        rom_memory[25631] = 3'b111;
        rom_memory[25632] = 3'b111;
        rom_memory[25633] = 3'b111;
        rom_memory[25634] = 3'b111;
        rom_memory[25635] = 3'b111;
        rom_memory[25636] = 3'b111;
        rom_memory[25637] = 3'b111;
        rom_memory[25638] = 3'b111;
        rom_memory[25639] = 3'b111;
        rom_memory[25640] = 3'b111;
        rom_memory[25641] = 3'b111;
        rom_memory[25642] = 3'b111;
        rom_memory[25643] = 3'b111;
        rom_memory[25644] = 3'b111;
        rom_memory[25645] = 3'b111;
        rom_memory[25646] = 3'b111;
        rom_memory[25647] = 3'b111;
        rom_memory[25648] = 3'b111;
        rom_memory[25649] = 3'b111;
        rom_memory[25650] = 3'b111;
        rom_memory[25651] = 3'b111;
        rom_memory[25652] = 3'b111;
        rom_memory[25653] = 3'b111;
        rom_memory[25654] = 3'b111;
        rom_memory[25655] = 3'b111;
        rom_memory[25656] = 3'b111;
        rom_memory[25657] = 3'b111;
        rom_memory[25658] = 3'b111;
        rom_memory[25659] = 3'b111;
        rom_memory[25660] = 3'b111;
        rom_memory[25661] = 3'b111;
        rom_memory[25662] = 3'b111;
        rom_memory[25663] = 3'b111;
        rom_memory[25664] = 3'b111;
        rom_memory[25665] = 3'b111;
        rom_memory[25666] = 3'b111;
        rom_memory[25667] = 3'b111;
        rom_memory[25668] = 3'b111;
        rom_memory[25669] = 3'b111;
        rom_memory[25670] = 3'b111;
        rom_memory[25671] = 3'b111;
        rom_memory[25672] = 3'b111;
        rom_memory[25673] = 3'b111;
        rom_memory[25674] = 3'b111;
        rom_memory[25675] = 3'b111;
        rom_memory[25676] = 3'b111;
        rom_memory[25677] = 3'b111;
        rom_memory[25678] = 3'b111;
        rom_memory[25679] = 3'b111;
        rom_memory[25680] = 3'b110;
        rom_memory[25681] = 3'b110;
        rom_memory[25682] = 3'b110;
        rom_memory[25683] = 3'b110;
        rom_memory[25684] = 3'b110;
        rom_memory[25685] = 3'b110;
        rom_memory[25686] = 3'b110;
        rom_memory[25687] = 3'b110;
        rom_memory[25688] = 3'b110;
        rom_memory[25689] = 3'b110;
        rom_memory[25690] = 3'b110;
        rom_memory[25691] = 3'b110;
        rom_memory[25692] = 3'b110;
        rom_memory[25693] = 3'b110;
        rom_memory[25694] = 3'b110;
        rom_memory[25695] = 3'b110;
        rom_memory[25696] = 3'b110;
        rom_memory[25697] = 3'b110;
        rom_memory[25698] = 3'b110;
        rom_memory[25699] = 3'b110;
        rom_memory[25700] = 3'b110;
        rom_memory[25701] = 3'b110;
        rom_memory[25702] = 3'b110;
        rom_memory[25703] = 3'b110;
        rom_memory[25704] = 3'b110;
        rom_memory[25705] = 3'b110;
        rom_memory[25706] = 3'b110;
        rom_memory[25707] = 3'b110;
        rom_memory[25708] = 3'b110;
        rom_memory[25709] = 3'b111;
        rom_memory[25710] = 3'b111;
        rom_memory[25711] = 3'b111;
        rom_memory[25712] = 3'b111;
        rom_memory[25713] = 3'b111;
        rom_memory[25714] = 3'b111;
        rom_memory[25715] = 3'b111;
        rom_memory[25716] = 3'b111;
        rom_memory[25717] = 3'b111;
        rom_memory[25718] = 3'b111;
        rom_memory[25719] = 3'b111;
        rom_memory[25720] = 3'b111;
        rom_memory[25721] = 3'b111;
        rom_memory[25722] = 3'b111;
        rom_memory[25723] = 3'b111;
        rom_memory[25724] = 3'b111;
        rom_memory[25725] = 3'b111;
        rom_memory[25726] = 3'b111;
        rom_memory[25727] = 3'b111;
        rom_memory[25728] = 3'b111;
        rom_memory[25729] = 3'b111;
        rom_memory[25730] = 3'b111;
        rom_memory[25731] = 3'b111;
        rom_memory[25732] = 3'b111;
        rom_memory[25733] = 3'b111;
        rom_memory[25734] = 3'b111;
        rom_memory[25735] = 3'b110;
        rom_memory[25736] = 3'b110;
        rom_memory[25737] = 3'b110;
        rom_memory[25738] = 3'b110;
        rom_memory[25739] = 3'b110;
        rom_memory[25740] = 3'b110;
        rom_memory[25741] = 3'b110;
        rom_memory[25742] = 3'b100;
        rom_memory[25743] = 3'b100;
        rom_memory[25744] = 3'b100;
        rom_memory[25745] = 3'b100;
        rom_memory[25746] = 3'b100;
        rom_memory[25747] = 3'b100;
        rom_memory[25748] = 3'b110;
        rom_memory[25749] = 3'b110;
        rom_memory[25750] = 3'b110;
        rom_memory[25751] = 3'b110;
        rom_memory[25752] = 3'b110;
        rom_memory[25753] = 3'b110;
        rom_memory[25754] = 3'b110;
        rom_memory[25755] = 3'b110;
        rom_memory[25756] = 3'b110;
        rom_memory[25757] = 3'b110;
        rom_memory[25758] = 3'b110;
        rom_memory[25759] = 3'b110;
        rom_memory[25760] = 3'b110;
        rom_memory[25761] = 3'b110;
        rom_memory[25762] = 3'b110;
        rom_memory[25763] = 3'b110;
        rom_memory[25764] = 3'b110;
        rom_memory[25765] = 3'b110;
        rom_memory[25766] = 3'b110;
        rom_memory[25767] = 3'b110;
        rom_memory[25768] = 3'b110;
        rom_memory[25769] = 3'b110;
        rom_memory[25770] = 3'b110;
        rom_memory[25771] = 3'b110;
        rom_memory[25772] = 3'b110;
        rom_memory[25773] = 3'b110;
        rom_memory[25774] = 3'b110;
        rom_memory[25775] = 3'b110;
        rom_memory[25776] = 3'b110;
        rom_memory[25777] = 3'b110;
        rom_memory[25778] = 3'b110;
        rom_memory[25779] = 3'b110;
        rom_memory[25780] = 3'b110;
        rom_memory[25781] = 3'b110;
        rom_memory[25782] = 3'b110;
        rom_memory[25783] = 3'b110;
        rom_memory[25784] = 3'b110;
        rom_memory[25785] = 3'b110;
        rom_memory[25786] = 3'b110;
        rom_memory[25787] = 3'b110;
        rom_memory[25788] = 3'b110;
        rom_memory[25789] = 3'b110;
        rom_memory[25790] = 3'b110;
        rom_memory[25791] = 3'b110;
        rom_memory[25792] = 3'b110;
        rom_memory[25793] = 3'b110;
        rom_memory[25794] = 3'b110;
        rom_memory[25795] = 3'b110;
        rom_memory[25796] = 3'b110;
        rom_memory[25797] = 3'b111;
        rom_memory[25798] = 3'b111;
        rom_memory[25799] = 3'b110;
        rom_memory[25800] = 3'b100;
        rom_memory[25801] = 3'b000;
        rom_memory[25802] = 3'b000;
        rom_memory[25803] = 3'b000;
        rom_memory[25804] = 3'b000;
        rom_memory[25805] = 3'b000;
        rom_memory[25806] = 3'b000;
        rom_memory[25807] = 3'b000;
        rom_memory[25808] = 3'b000;
        rom_memory[25809] = 3'b000;
        rom_memory[25810] = 3'b000;
        rom_memory[25811] = 3'b000;
        rom_memory[25812] = 3'b111;
        rom_memory[25813] = 3'b110;
        rom_memory[25814] = 3'b110;
        rom_memory[25815] = 3'b110;
        rom_memory[25816] = 3'b110;
        rom_memory[25817] = 3'b110;
        rom_memory[25818] = 3'b110;
        rom_memory[25819] = 3'b110;
        rom_memory[25820] = 3'b110;
        rom_memory[25821] = 3'b110;
        rom_memory[25822] = 3'b110;
        rom_memory[25823] = 3'b110;
        rom_memory[25824] = 3'b110;
        rom_memory[25825] = 3'b110;
        rom_memory[25826] = 3'b110;
        rom_memory[25827] = 3'b110;
        rom_memory[25828] = 3'b110;
        rom_memory[25829] = 3'b110;
        rom_memory[25830] = 3'b110;
        rom_memory[25831] = 3'b110;
        rom_memory[25832] = 3'b110;
        rom_memory[25833] = 3'b110;
        rom_memory[25834] = 3'b110;
        rom_memory[25835] = 3'b110;
        rom_memory[25836] = 3'b110;
        rom_memory[25837] = 3'b110;
        rom_memory[25838] = 3'b110;
        rom_memory[25839] = 3'b110;
        rom_memory[25840] = 3'b110;
        rom_memory[25841] = 3'b110;
        rom_memory[25842] = 3'b110;
        rom_memory[25843] = 3'b110;
        rom_memory[25844] = 3'b110;
        rom_memory[25845] = 3'b110;
        rom_memory[25846] = 3'b110;
        rom_memory[25847] = 3'b110;
        rom_memory[25848] = 3'b110;
        rom_memory[25849] = 3'b111;
        rom_memory[25850] = 3'b111;
        rom_memory[25851] = 3'b111;
        rom_memory[25852] = 3'b111;
        rom_memory[25853] = 3'b111;
        rom_memory[25854] = 3'b111;
        rom_memory[25855] = 3'b111;
        rom_memory[25856] = 3'b111;
        rom_memory[25857] = 3'b111;
        rom_memory[25858] = 3'b111;
        rom_memory[25859] = 3'b111;
        rom_memory[25860] = 3'b111;
        rom_memory[25861] = 3'b111;
        rom_memory[25862] = 3'b110;
        rom_memory[25863] = 3'b111;
        rom_memory[25864] = 3'b111;
        rom_memory[25865] = 3'b111;
        rom_memory[25866] = 3'b111;
        rom_memory[25867] = 3'b111;
        rom_memory[25868] = 3'b111;
        rom_memory[25869] = 3'b111;
        rom_memory[25870] = 3'b111;
        rom_memory[25871] = 3'b111;
        rom_memory[25872] = 3'b111;
        rom_memory[25873] = 3'b111;
        rom_memory[25874] = 3'b111;
        rom_memory[25875] = 3'b111;
        rom_memory[25876] = 3'b111;
        rom_memory[25877] = 3'b111;
        rom_memory[25878] = 3'b111;
        rom_memory[25879] = 3'b111;
        rom_memory[25880] = 3'b111;
        rom_memory[25881] = 3'b111;
        rom_memory[25882] = 3'b111;
        rom_memory[25883] = 3'b111;
        rom_memory[25884] = 3'b111;
        rom_memory[25885] = 3'b111;
        rom_memory[25886] = 3'b111;
        rom_memory[25887] = 3'b111;
        rom_memory[25888] = 3'b111;
        rom_memory[25889] = 3'b111;
        rom_memory[25890] = 3'b111;
        rom_memory[25891] = 3'b111;
        rom_memory[25892] = 3'b111;
        rom_memory[25893] = 3'b111;
        rom_memory[25894] = 3'b111;
        rom_memory[25895] = 3'b111;
        rom_memory[25896] = 3'b111;
        rom_memory[25897] = 3'b111;
        rom_memory[25898] = 3'b111;
        rom_memory[25899] = 3'b111;
        rom_memory[25900] = 3'b111;
        rom_memory[25901] = 3'b111;
        rom_memory[25902] = 3'b111;
        rom_memory[25903] = 3'b111;
        rom_memory[25904] = 3'b111;
        rom_memory[25905] = 3'b111;
        rom_memory[25906] = 3'b111;
        rom_memory[25907] = 3'b111;
        rom_memory[25908] = 3'b111;
        rom_memory[25909] = 3'b111;
        rom_memory[25910] = 3'b111;
        rom_memory[25911] = 3'b111;
        rom_memory[25912] = 3'b111;
        rom_memory[25913] = 3'b111;
        rom_memory[25914] = 3'b111;
        rom_memory[25915] = 3'b111;
        rom_memory[25916] = 3'b111;
        rom_memory[25917] = 3'b111;
        rom_memory[25918] = 3'b111;
        rom_memory[25919] = 3'b111;
        rom_memory[25920] = 3'b110;
        rom_memory[25921] = 3'b110;
        rom_memory[25922] = 3'b110;
        rom_memory[25923] = 3'b110;
        rom_memory[25924] = 3'b110;
        rom_memory[25925] = 3'b110;
        rom_memory[25926] = 3'b110;
        rom_memory[25927] = 3'b110;
        rom_memory[25928] = 3'b110;
        rom_memory[25929] = 3'b110;
        rom_memory[25930] = 3'b110;
        rom_memory[25931] = 3'b110;
        rom_memory[25932] = 3'b110;
        rom_memory[25933] = 3'b110;
        rom_memory[25934] = 3'b110;
        rom_memory[25935] = 3'b110;
        rom_memory[25936] = 3'b110;
        rom_memory[25937] = 3'b110;
        rom_memory[25938] = 3'b110;
        rom_memory[25939] = 3'b110;
        rom_memory[25940] = 3'b110;
        rom_memory[25941] = 3'b110;
        rom_memory[25942] = 3'b110;
        rom_memory[25943] = 3'b110;
        rom_memory[25944] = 3'b110;
        rom_memory[25945] = 3'b110;
        rom_memory[25946] = 3'b110;
        rom_memory[25947] = 3'b110;
        rom_memory[25948] = 3'b110;
        rom_memory[25949] = 3'b111;
        rom_memory[25950] = 3'b111;
        rom_memory[25951] = 3'b111;
        rom_memory[25952] = 3'b111;
        rom_memory[25953] = 3'b111;
        rom_memory[25954] = 3'b111;
        rom_memory[25955] = 3'b111;
        rom_memory[25956] = 3'b111;
        rom_memory[25957] = 3'b111;
        rom_memory[25958] = 3'b111;
        rom_memory[25959] = 3'b111;
        rom_memory[25960] = 3'b111;
        rom_memory[25961] = 3'b111;
        rom_memory[25962] = 3'b111;
        rom_memory[25963] = 3'b111;
        rom_memory[25964] = 3'b111;
        rom_memory[25965] = 3'b111;
        rom_memory[25966] = 3'b111;
        rom_memory[25967] = 3'b111;
        rom_memory[25968] = 3'b111;
        rom_memory[25969] = 3'b111;
        rom_memory[25970] = 3'b111;
        rom_memory[25971] = 3'b111;
        rom_memory[25972] = 3'b111;
        rom_memory[25973] = 3'b111;
        rom_memory[25974] = 3'b111;
        rom_memory[25975] = 3'b111;
        rom_memory[25976] = 3'b110;
        rom_memory[25977] = 3'b110;
        rom_memory[25978] = 3'b110;
        rom_memory[25979] = 3'b110;
        rom_memory[25980] = 3'b110;
        rom_memory[25981] = 3'b110;
        rom_memory[25982] = 3'b100;
        rom_memory[25983] = 3'b100;
        rom_memory[25984] = 3'b100;
        rom_memory[25985] = 3'b100;
        rom_memory[25986] = 3'b100;
        rom_memory[25987] = 3'b100;
        rom_memory[25988] = 3'b100;
        rom_memory[25989] = 3'b110;
        rom_memory[25990] = 3'b110;
        rom_memory[25991] = 3'b110;
        rom_memory[25992] = 3'b110;
        rom_memory[25993] = 3'b110;
        rom_memory[25994] = 3'b110;
        rom_memory[25995] = 3'b110;
        rom_memory[25996] = 3'b110;
        rom_memory[25997] = 3'b110;
        rom_memory[25998] = 3'b110;
        rom_memory[25999] = 3'b110;
        rom_memory[26000] = 3'b110;
        rom_memory[26001] = 3'b110;
        rom_memory[26002] = 3'b110;
        rom_memory[26003] = 3'b110;
        rom_memory[26004] = 3'b110;
        rom_memory[26005] = 3'b110;
        rom_memory[26006] = 3'b110;
        rom_memory[26007] = 3'b110;
        rom_memory[26008] = 3'b110;
        rom_memory[26009] = 3'b110;
        rom_memory[26010] = 3'b110;
        rom_memory[26011] = 3'b110;
        rom_memory[26012] = 3'b110;
        rom_memory[26013] = 3'b110;
        rom_memory[26014] = 3'b110;
        rom_memory[26015] = 3'b110;
        rom_memory[26016] = 3'b110;
        rom_memory[26017] = 3'b110;
        rom_memory[26018] = 3'b110;
        rom_memory[26019] = 3'b110;
        rom_memory[26020] = 3'b110;
        rom_memory[26021] = 3'b110;
        rom_memory[26022] = 3'b100;
        rom_memory[26023] = 3'b110;
        rom_memory[26024] = 3'b110;
        rom_memory[26025] = 3'b110;
        rom_memory[26026] = 3'b110;
        rom_memory[26027] = 3'b110;
        rom_memory[26028] = 3'b110;
        rom_memory[26029] = 3'b110;
        rom_memory[26030] = 3'b110;
        rom_memory[26031] = 3'b110;
        rom_memory[26032] = 3'b110;
        rom_memory[26033] = 3'b110;
        rom_memory[26034] = 3'b110;
        rom_memory[26035] = 3'b110;
        rom_memory[26036] = 3'b110;
        rom_memory[26037] = 3'b110;
        rom_memory[26038] = 3'b111;
        rom_memory[26039] = 3'b110;
        rom_memory[26040] = 3'b110;
        rom_memory[26041] = 3'b000;
        rom_memory[26042] = 3'b000;
        rom_memory[26043] = 3'b000;
        rom_memory[26044] = 3'b000;
        rom_memory[26045] = 3'b000;
        rom_memory[26046] = 3'b000;
        rom_memory[26047] = 3'b000;
        rom_memory[26048] = 3'b000;
        rom_memory[26049] = 3'b000;
        rom_memory[26050] = 3'b000;
        rom_memory[26051] = 3'b000;
        rom_memory[26052] = 3'b110;
        rom_memory[26053] = 3'b110;
        rom_memory[26054] = 3'b110;
        rom_memory[26055] = 3'b110;
        rom_memory[26056] = 3'b110;
        rom_memory[26057] = 3'b110;
        rom_memory[26058] = 3'b110;
        rom_memory[26059] = 3'b110;
        rom_memory[26060] = 3'b110;
        rom_memory[26061] = 3'b110;
        rom_memory[26062] = 3'b110;
        rom_memory[26063] = 3'b110;
        rom_memory[26064] = 3'b110;
        rom_memory[26065] = 3'b110;
        rom_memory[26066] = 3'b110;
        rom_memory[26067] = 3'b110;
        rom_memory[26068] = 3'b110;
        rom_memory[26069] = 3'b110;
        rom_memory[26070] = 3'b110;
        rom_memory[26071] = 3'b110;
        rom_memory[26072] = 3'b110;
        rom_memory[26073] = 3'b110;
        rom_memory[26074] = 3'b110;
        rom_memory[26075] = 3'b110;
        rom_memory[26076] = 3'b110;
        rom_memory[26077] = 3'b110;
        rom_memory[26078] = 3'b110;
        rom_memory[26079] = 3'b110;
        rom_memory[26080] = 3'b110;
        rom_memory[26081] = 3'b110;
        rom_memory[26082] = 3'b110;
        rom_memory[26083] = 3'b110;
        rom_memory[26084] = 3'b110;
        rom_memory[26085] = 3'b110;
        rom_memory[26086] = 3'b110;
        rom_memory[26087] = 3'b110;
        rom_memory[26088] = 3'b110;
        rom_memory[26089] = 3'b110;
        rom_memory[26090] = 3'b110;
        rom_memory[26091] = 3'b111;
        rom_memory[26092] = 3'b111;
        rom_memory[26093] = 3'b111;
        rom_memory[26094] = 3'b110;
        rom_memory[26095] = 3'b111;
        rom_memory[26096] = 3'b111;
        rom_memory[26097] = 3'b111;
        rom_memory[26098] = 3'b111;
        rom_memory[26099] = 3'b111;
        rom_memory[26100] = 3'b111;
        rom_memory[26101] = 3'b111;
        rom_memory[26102] = 3'b110;
        rom_memory[26103] = 3'b111;
        rom_memory[26104] = 3'b111;
        rom_memory[26105] = 3'b111;
        rom_memory[26106] = 3'b111;
        rom_memory[26107] = 3'b111;
        rom_memory[26108] = 3'b111;
        rom_memory[26109] = 3'b111;
        rom_memory[26110] = 3'b111;
        rom_memory[26111] = 3'b111;
        rom_memory[26112] = 3'b111;
        rom_memory[26113] = 3'b111;
        rom_memory[26114] = 3'b111;
        rom_memory[26115] = 3'b111;
        rom_memory[26116] = 3'b111;
        rom_memory[26117] = 3'b111;
        rom_memory[26118] = 3'b111;
        rom_memory[26119] = 3'b111;
        rom_memory[26120] = 3'b111;
        rom_memory[26121] = 3'b111;
        rom_memory[26122] = 3'b111;
        rom_memory[26123] = 3'b111;
        rom_memory[26124] = 3'b111;
        rom_memory[26125] = 3'b111;
        rom_memory[26126] = 3'b111;
        rom_memory[26127] = 3'b111;
        rom_memory[26128] = 3'b111;
        rom_memory[26129] = 3'b111;
        rom_memory[26130] = 3'b111;
        rom_memory[26131] = 3'b111;
        rom_memory[26132] = 3'b111;
        rom_memory[26133] = 3'b111;
        rom_memory[26134] = 3'b111;
        rom_memory[26135] = 3'b111;
        rom_memory[26136] = 3'b111;
        rom_memory[26137] = 3'b111;
        rom_memory[26138] = 3'b111;
        rom_memory[26139] = 3'b111;
        rom_memory[26140] = 3'b111;
        rom_memory[26141] = 3'b111;
        rom_memory[26142] = 3'b111;
        rom_memory[26143] = 3'b111;
        rom_memory[26144] = 3'b111;
        rom_memory[26145] = 3'b111;
        rom_memory[26146] = 3'b111;
        rom_memory[26147] = 3'b111;
        rom_memory[26148] = 3'b111;
        rom_memory[26149] = 3'b111;
        rom_memory[26150] = 3'b111;
        rom_memory[26151] = 3'b111;
        rom_memory[26152] = 3'b111;
        rom_memory[26153] = 3'b111;
        rom_memory[26154] = 3'b111;
        rom_memory[26155] = 3'b111;
        rom_memory[26156] = 3'b111;
        rom_memory[26157] = 3'b111;
        rom_memory[26158] = 3'b111;
        rom_memory[26159] = 3'b111;
        rom_memory[26160] = 3'b110;
        rom_memory[26161] = 3'b110;
        rom_memory[26162] = 3'b110;
        rom_memory[26163] = 3'b110;
        rom_memory[26164] = 3'b110;
        rom_memory[26165] = 3'b110;
        rom_memory[26166] = 3'b110;
        rom_memory[26167] = 3'b110;
        rom_memory[26168] = 3'b110;
        rom_memory[26169] = 3'b110;
        rom_memory[26170] = 3'b110;
        rom_memory[26171] = 3'b110;
        rom_memory[26172] = 3'b110;
        rom_memory[26173] = 3'b110;
        rom_memory[26174] = 3'b110;
        rom_memory[26175] = 3'b110;
        rom_memory[26176] = 3'b110;
        rom_memory[26177] = 3'b110;
        rom_memory[26178] = 3'b110;
        rom_memory[26179] = 3'b110;
        rom_memory[26180] = 3'b110;
        rom_memory[26181] = 3'b110;
        rom_memory[26182] = 3'b110;
        rom_memory[26183] = 3'b110;
        rom_memory[26184] = 3'b110;
        rom_memory[26185] = 3'b110;
        rom_memory[26186] = 3'b110;
        rom_memory[26187] = 3'b110;
        rom_memory[26188] = 3'b110;
        rom_memory[26189] = 3'b110;
        rom_memory[26190] = 3'b111;
        rom_memory[26191] = 3'b111;
        rom_memory[26192] = 3'b111;
        rom_memory[26193] = 3'b111;
        rom_memory[26194] = 3'b111;
        rom_memory[26195] = 3'b111;
        rom_memory[26196] = 3'b111;
        rom_memory[26197] = 3'b111;
        rom_memory[26198] = 3'b111;
        rom_memory[26199] = 3'b111;
        rom_memory[26200] = 3'b111;
        rom_memory[26201] = 3'b111;
        rom_memory[26202] = 3'b111;
        rom_memory[26203] = 3'b111;
        rom_memory[26204] = 3'b111;
        rom_memory[26205] = 3'b111;
        rom_memory[26206] = 3'b111;
        rom_memory[26207] = 3'b111;
        rom_memory[26208] = 3'b111;
        rom_memory[26209] = 3'b111;
        rom_memory[26210] = 3'b111;
        rom_memory[26211] = 3'b111;
        rom_memory[26212] = 3'b111;
        rom_memory[26213] = 3'b111;
        rom_memory[26214] = 3'b111;
        rom_memory[26215] = 3'b111;
        rom_memory[26216] = 3'b110;
        rom_memory[26217] = 3'b110;
        rom_memory[26218] = 3'b110;
        rom_memory[26219] = 3'b110;
        rom_memory[26220] = 3'b110;
        rom_memory[26221] = 3'b110;
        rom_memory[26222] = 3'b110;
        rom_memory[26223] = 3'b110;
        rom_memory[26224] = 3'b100;
        rom_memory[26225] = 3'b100;
        rom_memory[26226] = 3'b100;
        rom_memory[26227] = 3'b100;
        rom_memory[26228] = 3'b110;
        rom_memory[26229] = 3'b110;
        rom_memory[26230] = 3'b110;
        rom_memory[26231] = 3'b110;
        rom_memory[26232] = 3'b110;
        rom_memory[26233] = 3'b110;
        rom_memory[26234] = 3'b110;
        rom_memory[26235] = 3'b110;
        rom_memory[26236] = 3'b110;
        rom_memory[26237] = 3'b110;
        rom_memory[26238] = 3'b110;
        rom_memory[26239] = 3'b110;
        rom_memory[26240] = 3'b110;
        rom_memory[26241] = 3'b110;
        rom_memory[26242] = 3'b110;
        rom_memory[26243] = 3'b110;
        rom_memory[26244] = 3'b110;
        rom_memory[26245] = 3'b110;
        rom_memory[26246] = 3'b110;
        rom_memory[26247] = 3'b110;
        rom_memory[26248] = 3'b110;
        rom_memory[26249] = 3'b110;
        rom_memory[26250] = 3'b110;
        rom_memory[26251] = 3'b110;
        rom_memory[26252] = 3'b110;
        rom_memory[26253] = 3'b110;
        rom_memory[26254] = 3'b110;
        rom_memory[26255] = 3'b110;
        rom_memory[26256] = 3'b110;
        rom_memory[26257] = 3'b110;
        rom_memory[26258] = 3'b110;
        rom_memory[26259] = 3'b110;
        rom_memory[26260] = 3'b110;
        rom_memory[26261] = 3'b110;
        rom_memory[26262] = 3'b110;
        rom_memory[26263] = 3'b110;
        rom_memory[26264] = 3'b110;
        rom_memory[26265] = 3'b110;
        rom_memory[26266] = 3'b110;
        rom_memory[26267] = 3'b110;
        rom_memory[26268] = 3'b110;
        rom_memory[26269] = 3'b110;
        rom_memory[26270] = 3'b110;
        rom_memory[26271] = 3'b110;
        rom_memory[26272] = 3'b110;
        rom_memory[26273] = 3'b110;
        rom_memory[26274] = 3'b110;
        rom_memory[26275] = 3'b110;
        rom_memory[26276] = 3'b110;
        rom_memory[26277] = 3'b110;
        rom_memory[26278] = 3'b110;
        rom_memory[26279] = 3'b110;
        rom_memory[26280] = 3'b110;
        rom_memory[26281] = 3'b110;
        rom_memory[26282] = 3'b000;
        rom_memory[26283] = 3'b000;
        rom_memory[26284] = 3'b000;
        rom_memory[26285] = 3'b000;
        rom_memory[26286] = 3'b000;
        rom_memory[26287] = 3'b000;
        rom_memory[26288] = 3'b000;
        rom_memory[26289] = 3'b000;
        rom_memory[26290] = 3'b000;
        rom_memory[26291] = 3'b000;
        rom_memory[26292] = 3'b100;
        rom_memory[26293] = 3'b110;
        rom_memory[26294] = 3'b110;
        rom_memory[26295] = 3'b110;
        rom_memory[26296] = 3'b110;
        rom_memory[26297] = 3'b110;
        rom_memory[26298] = 3'b110;
        rom_memory[26299] = 3'b110;
        rom_memory[26300] = 3'b110;
        rom_memory[26301] = 3'b110;
        rom_memory[26302] = 3'b110;
        rom_memory[26303] = 3'b110;
        rom_memory[26304] = 3'b110;
        rom_memory[26305] = 3'b110;
        rom_memory[26306] = 3'b110;
        rom_memory[26307] = 3'b110;
        rom_memory[26308] = 3'b110;
        rom_memory[26309] = 3'b110;
        rom_memory[26310] = 3'b110;
        rom_memory[26311] = 3'b110;
        rom_memory[26312] = 3'b110;
        rom_memory[26313] = 3'b110;
        rom_memory[26314] = 3'b110;
        rom_memory[26315] = 3'b110;
        rom_memory[26316] = 3'b110;
        rom_memory[26317] = 3'b110;
        rom_memory[26318] = 3'b110;
        rom_memory[26319] = 3'b110;
        rom_memory[26320] = 3'b110;
        rom_memory[26321] = 3'b110;
        rom_memory[26322] = 3'b110;
        rom_memory[26323] = 3'b110;
        rom_memory[26324] = 3'b110;
        rom_memory[26325] = 3'b110;
        rom_memory[26326] = 3'b110;
        rom_memory[26327] = 3'b110;
        rom_memory[26328] = 3'b110;
        rom_memory[26329] = 3'b110;
        rom_memory[26330] = 3'b110;
        rom_memory[26331] = 3'b111;
        rom_memory[26332] = 3'b111;
        rom_memory[26333] = 3'b111;
        rom_memory[26334] = 3'b110;
        rom_memory[26335] = 3'b110;
        rom_memory[26336] = 3'b110;
        rom_memory[26337] = 3'b111;
        rom_memory[26338] = 3'b111;
        rom_memory[26339] = 3'b111;
        rom_memory[26340] = 3'b111;
        rom_memory[26341] = 3'b111;
        rom_memory[26342] = 3'b111;
        rom_memory[26343] = 3'b111;
        rom_memory[26344] = 3'b111;
        rom_memory[26345] = 3'b111;
        rom_memory[26346] = 3'b111;
        rom_memory[26347] = 3'b111;
        rom_memory[26348] = 3'b111;
        rom_memory[26349] = 3'b111;
        rom_memory[26350] = 3'b111;
        rom_memory[26351] = 3'b111;
        rom_memory[26352] = 3'b111;
        rom_memory[26353] = 3'b111;
        rom_memory[26354] = 3'b111;
        rom_memory[26355] = 3'b111;
        rom_memory[26356] = 3'b111;
        rom_memory[26357] = 3'b111;
        rom_memory[26358] = 3'b111;
        rom_memory[26359] = 3'b111;
        rom_memory[26360] = 3'b111;
        rom_memory[26361] = 3'b111;
        rom_memory[26362] = 3'b111;
        rom_memory[26363] = 3'b111;
        rom_memory[26364] = 3'b111;
        rom_memory[26365] = 3'b111;
        rom_memory[26366] = 3'b111;
        rom_memory[26367] = 3'b111;
        rom_memory[26368] = 3'b111;
        rom_memory[26369] = 3'b111;
        rom_memory[26370] = 3'b111;
        rom_memory[26371] = 3'b111;
        rom_memory[26372] = 3'b111;
        rom_memory[26373] = 3'b111;
        rom_memory[26374] = 3'b111;
        rom_memory[26375] = 3'b111;
        rom_memory[26376] = 3'b111;
        rom_memory[26377] = 3'b111;
        rom_memory[26378] = 3'b111;
        rom_memory[26379] = 3'b111;
        rom_memory[26380] = 3'b111;
        rom_memory[26381] = 3'b111;
        rom_memory[26382] = 3'b111;
        rom_memory[26383] = 3'b111;
        rom_memory[26384] = 3'b111;
        rom_memory[26385] = 3'b111;
        rom_memory[26386] = 3'b111;
        rom_memory[26387] = 3'b111;
        rom_memory[26388] = 3'b111;
        rom_memory[26389] = 3'b111;
        rom_memory[26390] = 3'b111;
        rom_memory[26391] = 3'b111;
        rom_memory[26392] = 3'b111;
        rom_memory[26393] = 3'b111;
        rom_memory[26394] = 3'b111;
        rom_memory[26395] = 3'b111;
        rom_memory[26396] = 3'b111;
        rom_memory[26397] = 3'b111;
        rom_memory[26398] = 3'b111;
        rom_memory[26399] = 3'b111;
        rom_memory[26400] = 3'b110;
        rom_memory[26401] = 3'b110;
        rom_memory[26402] = 3'b110;
        rom_memory[26403] = 3'b110;
        rom_memory[26404] = 3'b110;
        rom_memory[26405] = 3'b110;
        rom_memory[26406] = 3'b110;
        rom_memory[26407] = 3'b110;
        rom_memory[26408] = 3'b110;
        rom_memory[26409] = 3'b110;
        rom_memory[26410] = 3'b110;
        rom_memory[26411] = 3'b110;
        rom_memory[26412] = 3'b110;
        rom_memory[26413] = 3'b110;
        rom_memory[26414] = 3'b110;
        rom_memory[26415] = 3'b110;
        rom_memory[26416] = 3'b110;
        rom_memory[26417] = 3'b110;
        rom_memory[26418] = 3'b110;
        rom_memory[26419] = 3'b110;
        rom_memory[26420] = 3'b110;
        rom_memory[26421] = 3'b110;
        rom_memory[26422] = 3'b110;
        rom_memory[26423] = 3'b110;
        rom_memory[26424] = 3'b110;
        rom_memory[26425] = 3'b110;
        rom_memory[26426] = 3'b110;
        rom_memory[26427] = 3'b110;
        rom_memory[26428] = 3'b110;
        rom_memory[26429] = 3'b110;
        rom_memory[26430] = 3'b111;
        rom_memory[26431] = 3'b111;
        rom_memory[26432] = 3'b111;
        rom_memory[26433] = 3'b111;
        rom_memory[26434] = 3'b111;
        rom_memory[26435] = 3'b111;
        rom_memory[26436] = 3'b111;
        rom_memory[26437] = 3'b111;
        rom_memory[26438] = 3'b111;
        rom_memory[26439] = 3'b111;
        rom_memory[26440] = 3'b111;
        rom_memory[26441] = 3'b111;
        rom_memory[26442] = 3'b111;
        rom_memory[26443] = 3'b111;
        rom_memory[26444] = 3'b111;
        rom_memory[26445] = 3'b111;
        rom_memory[26446] = 3'b111;
        rom_memory[26447] = 3'b111;
        rom_memory[26448] = 3'b111;
        rom_memory[26449] = 3'b111;
        rom_memory[26450] = 3'b111;
        rom_memory[26451] = 3'b111;
        rom_memory[26452] = 3'b111;
        rom_memory[26453] = 3'b111;
        rom_memory[26454] = 3'b111;
        rom_memory[26455] = 3'b111;
        rom_memory[26456] = 3'b111;
        rom_memory[26457] = 3'b110;
        rom_memory[26458] = 3'b110;
        rom_memory[26459] = 3'b110;
        rom_memory[26460] = 3'b100;
        rom_memory[26461] = 3'b110;
        rom_memory[26462] = 3'b110;
        rom_memory[26463] = 3'b110;
        rom_memory[26464] = 3'b110;
        rom_memory[26465] = 3'b110;
        rom_memory[26466] = 3'b100;
        rom_memory[26467] = 3'b100;
        rom_memory[26468] = 3'b100;
        rom_memory[26469] = 3'b100;
        rom_memory[26470] = 3'b110;
        rom_memory[26471] = 3'b110;
        rom_memory[26472] = 3'b110;
        rom_memory[26473] = 3'b110;
        rom_memory[26474] = 3'b110;
        rom_memory[26475] = 3'b110;
        rom_memory[26476] = 3'b110;
        rom_memory[26477] = 3'b110;
        rom_memory[26478] = 3'b110;
        rom_memory[26479] = 3'b110;
        rom_memory[26480] = 3'b110;
        rom_memory[26481] = 3'b110;
        rom_memory[26482] = 3'b110;
        rom_memory[26483] = 3'b110;
        rom_memory[26484] = 3'b110;
        rom_memory[26485] = 3'b110;
        rom_memory[26486] = 3'b110;
        rom_memory[26487] = 3'b110;
        rom_memory[26488] = 3'b110;
        rom_memory[26489] = 3'b110;
        rom_memory[26490] = 3'b110;
        rom_memory[26491] = 3'b110;
        rom_memory[26492] = 3'b110;
        rom_memory[26493] = 3'b110;
        rom_memory[26494] = 3'b110;
        rom_memory[26495] = 3'b110;
        rom_memory[26496] = 3'b110;
        rom_memory[26497] = 3'b110;
        rom_memory[26498] = 3'b110;
        rom_memory[26499] = 3'b110;
        rom_memory[26500] = 3'b110;
        rom_memory[26501] = 3'b110;
        rom_memory[26502] = 3'b110;
        rom_memory[26503] = 3'b100;
        rom_memory[26504] = 3'b110;
        rom_memory[26505] = 3'b110;
        rom_memory[26506] = 3'b110;
        rom_memory[26507] = 3'b110;
        rom_memory[26508] = 3'b110;
        rom_memory[26509] = 3'b110;
        rom_memory[26510] = 3'b110;
        rom_memory[26511] = 3'b110;
        rom_memory[26512] = 3'b110;
        rom_memory[26513] = 3'b110;
        rom_memory[26514] = 3'b110;
        rom_memory[26515] = 3'b110;
        rom_memory[26516] = 3'b110;
        rom_memory[26517] = 3'b110;
        rom_memory[26518] = 3'b110;
        rom_memory[26519] = 3'b110;
        rom_memory[26520] = 3'b110;
        rom_memory[26521] = 3'b110;
        rom_memory[26522] = 3'b100;
        rom_memory[26523] = 3'b000;
        rom_memory[26524] = 3'b000;
        rom_memory[26525] = 3'b000;
        rom_memory[26526] = 3'b000;
        rom_memory[26527] = 3'b000;
        rom_memory[26528] = 3'b000;
        rom_memory[26529] = 3'b000;
        rom_memory[26530] = 3'b000;
        rom_memory[26531] = 3'b000;
        rom_memory[26532] = 3'b000;
        rom_memory[26533] = 3'b110;
        rom_memory[26534] = 3'b110;
        rom_memory[26535] = 3'b110;
        rom_memory[26536] = 3'b110;
        rom_memory[26537] = 3'b110;
        rom_memory[26538] = 3'b110;
        rom_memory[26539] = 3'b110;
        rom_memory[26540] = 3'b110;
        rom_memory[26541] = 3'b110;
        rom_memory[26542] = 3'b110;
        rom_memory[26543] = 3'b110;
        rom_memory[26544] = 3'b110;
        rom_memory[26545] = 3'b110;
        rom_memory[26546] = 3'b110;
        rom_memory[26547] = 3'b110;
        rom_memory[26548] = 3'b110;
        rom_memory[26549] = 3'b110;
        rom_memory[26550] = 3'b110;
        rom_memory[26551] = 3'b110;
        rom_memory[26552] = 3'b110;
        rom_memory[26553] = 3'b110;
        rom_memory[26554] = 3'b110;
        rom_memory[26555] = 3'b110;
        rom_memory[26556] = 3'b110;
        rom_memory[26557] = 3'b110;
        rom_memory[26558] = 3'b110;
        rom_memory[26559] = 3'b110;
        rom_memory[26560] = 3'b110;
        rom_memory[26561] = 3'b110;
        rom_memory[26562] = 3'b110;
        rom_memory[26563] = 3'b110;
        rom_memory[26564] = 3'b110;
        rom_memory[26565] = 3'b110;
        rom_memory[26566] = 3'b110;
        rom_memory[26567] = 3'b111;
        rom_memory[26568] = 3'b110;
        rom_memory[26569] = 3'b110;
        rom_memory[26570] = 3'b110;
        rom_memory[26571] = 3'b110;
        rom_memory[26572] = 3'b111;
        rom_memory[26573] = 3'b110;
        rom_memory[26574] = 3'b110;
        rom_memory[26575] = 3'b110;
        rom_memory[26576] = 3'b110;
        rom_memory[26577] = 3'b110;
        rom_memory[26578] = 3'b110;
        rom_memory[26579] = 3'b110;
        rom_memory[26580] = 3'b110;
        rom_memory[26581] = 3'b111;
        rom_memory[26582] = 3'b111;
        rom_memory[26583] = 3'b111;
        rom_memory[26584] = 3'b111;
        rom_memory[26585] = 3'b111;
        rom_memory[26586] = 3'b111;
        rom_memory[26587] = 3'b111;
        rom_memory[26588] = 3'b111;
        rom_memory[26589] = 3'b111;
        rom_memory[26590] = 3'b111;
        rom_memory[26591] = 3'b111;
        rom_memory[26592] = 3'b111;
        rom_memory[26593] = 3'b111;
        rom_memory[26594] = 3'b111;
        rom_memory[26595] = 3'b111;
        rom_memory[26596] = 3'b111;
        rom_memory[26597] = 3'b111;
        rom_memory[26598] = 3'b111;
        rom_memory[26599] = 3'b111;
        rom_memory[26600] = 3'b111;
        rom_memory[26601] = 3'b111;
        rom_memory[26602] = 3'b111;
        rom_memory[26603] = 3'b111;
        rom_memory[26604] = 3'b111;
        rom_memory[26605] = 3'b111;
        rom_memory[26606] = 3'b111;
        rom_memory[26607] = 3'b111;
        rom_memory[26608] = 3'b111;
        rom_memory[26609] = 3'b111;
        rom_memory[26610] = 3'b111;
        rom_memory[26611] = 3'b111;
        rom_memory[26612] = 3'b111;
        rom_memory[26613] = 3'b111;
        rom_memory[26614] = 3'b111;
        rom_memory[26615] = 3'b111;
        rom_memory[26616] = 3'b111;
        rom_memory[26617] = 3'b111;
        rom_memory[26618] = 3'b111;
        rom_memory[26619] = 3'b111;
        rom_memory[26620] = 3'b111;
        rom_memory[26621] = 3'b111;
        rom_memory[26622] = 3'b111;
        rom_memory[26623] = 3'b111;
        rom_memory[26624] = 3'b111;
        rom_memory[26625] = 3'b111;
        rom_memory[26626] = 3'b111;
        rom_memory[26627] = 3'b111;
        rom_memory[26628] = 3'b111;
        rom_memory[26629] = 3'b111;
        rom_memory[26630] = 3'b111;
        rom_memory[26631] = 3'b111;
        rom_memory[26632] = 3'b111;
        rom_memory[26633] = 3'b111;
        rom_memory[26634] = 3'b111;
        rom_memory[26635] = 3'b111;
        rom_memory[26636] = 3'b111;
        rom_memory[26637] = 3'b111;
        rom_memory[26638] = 3'b111;
        rom_memory[26639] = 3'b111;
        rom_memory[26640] = 3'b110;
        rom_memory[26641] = 3'b110;
        rom_memory[26642] = 3'b110;
        rom_memory[26643] = 3'b110;
        rom_memory[26644] = 3'b110;
        rom_memory[26645] = 3'b110;
        rom_memory[26646] = 3'b110;
        rom_memory[26647] = 3'b110;
        rom_memory[26648] = 3'b110;
        rom_memory[26649] = 3'b110;
        rom_memory[26650] = 3'b110;
        rom_memory[26651] = 3'b110;
        rom_memory[26652] = 3'b110;
        rom_memory[26653] = 3'b110;
        rom_memory[26654] = 3'b110;
        rom_memory[26655] = 3'b110;
        rom_memory[26656] = 3'b110;
        rom_memory[26657] = 3'b110;
        rom_memory[26658] = 3'b110;
        rom_memory[26659] = 3'b110;
        rom_memory[26660] = 3'b110;
        rom_memory[26661] = 3'b110;
        rom_memory[26662] = 3'b110;
        rom_memory[26663] = 3'b110;
        rom_memory[26664] = 3'b110;
        rom_memory[26665] = 3'b110;
        rom_memory[26666] = 3'b110;
        rom_memory[26667] = 3'b110;
        rom_memory[26668] = 3'b110;
        rom_memory[26669] = 3'b110;
        rom_memory[26670] = 3'b110;
        rom_memory[26671] = 3'b111;
        rom_memory[26672] = 3'b111;
        rom_memory[26673] = 3'b111;
        rom_memory[26674] = 3'b111;
        rom_memory[26675] = 3'b111;
        rom_memory[26676] = 3'b111;
        rom_memory[26677] = 3'b111;
        rom_memory[26678] = 3'b111;
        rom_memory[26679] = 3'b111;
        rom_memory[26680] = 3'b111;
        rom_memory[26681] = 3'b111;
        rom_memory[26682] = 3'b111;
        rom_memory[26683] = 3'b111;
        rom_memory[26684] = 3'b111;
        rom_memory[26685] = 3'b111;
        rom_memory[26686] = 3'b111;
        rom_memory[26687] = 3'b111;
        rom_memory[26688] = 3'b111;
        rom_memory[26689] = 3'b111;
        rom_memory[26690] = 3'b111;
        rom_memory[26691] = 3'b111;
        rom_memory[26692] = 3'b111;
        rom_memory[26693] = 3'b111;
        rom_memory[26694] = 3'b111;
        rom_memory[26695] = 3'b111;
        rom_memory[26696] = 3'b111;
        rom_memory[26697] = 3'b111;
        rom_memory[26698] = 3'b110;
        rom_memory[26699] = 3'b110;
        rom_memory[26700] = 3'b100;
        rom_memory[26701] = 3'b110;
        rom_memory[26702] = 3'b110;
        rom_memory[26703] = 3'b110;
        rom_memory[26704] = 3'b110;
        rom_memory[26705] = 3'b110;
        rom_memory[26706] = 3'b110;
        rom_memory[26707] = 3'b100;
        rom_memory[26708] = 3'b100;
        rom_memory[26709] = 3'b100;
        rom_memory[26710] = 3'b110;
        rom_memory[26711] = 3'b110;
        rom_memory[26712] = 3'b110;
        rom_memory[26713] = 3'b110;
        rom_memory[26714] = 3'b110;
        rom_memory[26715] = 3'b110;
        rom_memory[26716] = 3'b110;
        rom_memory[26717] = 3'b110;
        rom_memory[26718] = 3'b110;
        rom_memory[26719] = 3'b110;
        rom_memory[26720] = 3'b110;
        rom_memory[26721] = 3'b110;
        rom_memory[26722] = 3'b110;
        rom_memory[26723] = 3'b110;
        rom_memory[26724] = 3'b110;
        rom_memory[26725] = 3'b110;
        rom_memory[26726] = 3'b110;
        rom_memory[26727] = 3'b110;
        rom_memory[26728] = 3'b110;
        rom_memory[26729] = 3'b110;
        rom_memory[26730] = 3'b110;
        rom_memory[26731] = 3'b110;
        rom_memory[26732] = 3'b110;
        rom_memory[26733] = 3'b110;
        rom_memory[26734] = 3'b110;
        rom_memory[26735] = 3'b110;
        rom_memory[26736] = 3'b110;
        rom_memory[26737] = 3'b110;
        rom_memory[26738] = 3'b110;
        rom_memory[26739] = 3'b110;
        rom_memory[26740] = 3'b110;
        rom_memory[26741] = 3'b110;
        rom_memory[26742] = 3'b110;
        rom_memory[26743] = 3'b110;
        rom_memory[26744] = 3'b110;
        rom_memory[26745] = 3'b110;
        rom_memory[26746] = 3'b110;
        rom_memory[26747] = 3'b110;
        rom_memory[26748] = 3'b110;
        rom_memory[26749] = 3'b110;
        rom_memory[26750] = 3'b110;
        rom_memory[26751] = 3'b110;
        rom_memory[26752] = 3'b110;
        rom_memory[26753] = 3'b110;
        rom_memory[26754] = 3'b110;
        rom_memory[26755] = 3'b110;
        rom_memory[26756] = 3'b110;
        rom_memory[26757] = 3'b110;
        rom_memory[26758] = 3'b110;
        rom_memory[26759] = 3'b110;
        rom_memory[26760] = 3'b110;
        rom_memory[26761] = 3'b110;
        rom_memory[26762] = 3'b100;
        rom_memory[26763] = 3'b000;
        rom_memory[26764] = 3'b100;
        rom_memory[26765] = 3'b100;
        rom_memory[26766] = 3'b000;
        rom_memory[26767] = 3'b000;
        rom_memory[26768] = 3'b000;
        rom_memory[26769] = 3'b000;
        rom_memory[26770] = 3'b000;
        rom_memory[26771] = 3'b000;
        rom_memory[26772] = 3'b000;
        rom_memory[26773] = 3'b110;
        rom_memory[26774] = 3'b110;
        rom_memory[26775] = 3'b110;
        rom_memory[26776] = 3'b110;
        rom_memory[26777] = 3'b110;
        rom_memory[26778] = 3'b110;
        rom_memory[26779] = 3'b110;
        rom_memory[26780] = 3'b110;
        rom_memory[26781] = 3'b110;
        rom_memory[26782] = 3'b110;
        rom_memory[26783] = 3'b110;
        rom_memory[26784] = 3'b110;
        rom_memory[26785] = 3'b110;
        rom_memory[26786] = 3'b110;
        rom_memory[26787] = 3'b110;
        rom_memory[26788] = 3'b110;
        rom_memory[26789] = 3'b110;
        rom_memory[26790] = 3'b110;
        rom_memory[26791] = 3'b110;
        rom_memory[26792] = 3'b110;
        rom_memory[26793] = 3'b110;
        rom_memory[26794] = 3'b110;
        rom_memory[26795] = 3'b110;
        rom_memory[26796] = 3'b110;
        rom_memory[26797] = 3'b110;
        rom_memory[26798] = 3'b110;
        rom_memory[26799] = 3'b110;
        rom_memory[26800] = 3'b110;
        rom_memory[26801] = 3'b110;
        rom_memory[26802] = 3'b110;
        rom_memory[26803] = 3'b110;
        rom_memory[26804] = 3'b110;
        rom_memory[26805] = 3'b110;
        rom_memory[26806] = 3'b110;
        rom_memory[26807] = 3'b110;
        rom_memory[26808] = 3'b110;
        rom_memory[26809] = 3'b110;
        rom_memory[26810] = 3'b110;
        rom_memory[26811] = 3'b111;
        rom_memory[26812] = 3'b110;
        rom_memory[26813] = 3'b110;
        rom_memory[26814] = 3'b110;
        rom_memory[26815] = 3'b110;
        rom_memory[26816] = 3'b110;
        rom_memory[26817] = 3'b110;
        rom_memory[26818] = 3'b111;
        rom_memory[26819] = 3'b111;
        rom_memory[26820] = 3'b110;
        rom_memory[26821] = 3'b110;
        rom_memory[26822] = 3'b111;
        rom_memory[26823] = 3'b111;
        rom_memory[26824] = 3'b111;
        rom_memory[26825] = 3'b111;
        rom_memory[26826] = 3'b111;
        rom_memory[26827] = 3'b111;
        rom_memory[26828] = 3'b111;
        rom_memory[26829] = 3'b111;
        rom_memory[26830] = 3'b111;
        rom_memory[26831] = 3'b111;
        rom_memory[26832] = 3'b111;
        rom_memory[26833] = 3'b111;
        rom_memory[26834] = 3'b111;
        rom_memory[26835] = 3'b111;
        rom_memory[26836] = 3'b111;
        rom_memory[26837] = 3'b111;
        rom_memory[26838] = 3'b111;
        rom_memory[26839] = 3'b111;
        rom_memory[26840] = 3'b111;
        rom_memory[26841] = 3'b111;
        rom_memory[26842] = 3'b111;
        rom_memory[26843] = 3'b111;
        rom_memory[26844] = 3'b111;
        rom_memory[26845] = 3'b111;
        rom_memory[26846] = 3'b111;
        rom_memory[26847] = 3'b111;
        rom_memory[26848] = 3'b111;
        rom_memory[26849] = 3'b111;
        rom_memory[26850] = 3'b111;
        rom_memory[26851] = 3'b111;
        rom_memory[26852] = 3'b111;
        rom_memory[26853] = 3'b111;
        rom_memory[26854] = 3'b111;
        rom_memory[26855] = 3'b111;
        rom_memory[26856] = 3'b111;
        rom_memory[26857] = 3'b111;
        rom_memory[26858] = 3'b111;
        rom_memory[26859] = 3'b111;
        rom_memory[26860] = 3'b111;
        rom_memory[26861] = 3'b111;
        rom_memory[26862] = 3'b111;
        rom_memory[26863] = 3'b111;
        rom_memory[26864] = 3'b111;
        rom_memory[26865] = 3'b111;
        rom_memory[26866] = 3'b111;
        rom_memory[26867] = 3'b111;
        rom_memory[26868] = 3'b111;
        rom_memory[26869] = 3'b111;
        rom_memory[26870] = 3'b111;
        rom_memory[26871] = 3'b111;
        rom_memory[26872] = 3'b111;
        rom_memory[26873] = 3'b111;
        rom_memory[26874] = 3'b111;
        rom_memory[26875] = 3'b111;
        rom_memory[26876] = 3'b111;
        rom_memory[26877] = 3'b111;
        rom_memory[26878] = 3'b111;
        rom_memory[26879] = 3'b111;
        rom_memory[26880] = 3'b110;
        rom_memory[26881] = 3'b110;
        rom_memory[26882] = 3'b110;
        rom_memory[26883] = 3'b110;
        rom_memory[26884] = 3'b110;
        rom_memory[26885] = 3'b110;
        rom_memory[26886] = 3'b110;
        rom_memory[26887] = 3'b110;
        rom_memory[26888] = 3'b110;
        rom_memory[26889] = 3'b110;
        rom_memory[26890] = 3'b110;
        rom_memory[26891] = 3'b110;
        rom_memory[26892] = 3'b110;
        rom_memory[26893] = 3'b110;
        rom_memory[26894] = 3'b110;
        rom_memory[26895] = 3'b110;
        rom_memory[26896] = 3'b110;
        rom_memory[26897] = 3'b110;
        rom_memory[26898] = 3'b110;
        rom_memory[26899] = 3'b110;
        rom_memory[26900] = 3'b110;
        rom_memory[26901] = 3'b110;
        rom_memory[26902] = 3'b110;
        rom_memory[26903] = 3'b110;
        rom_memory[26904] = 3'b110;
        rom_memory[26905] = 3'b110;
        rom_memory[26906] = 3'b110;
        rom_memory[26907] = 3'b110;
        rom_memory[26908] = 3'b110;
        rom_memory[26909] = 3'b110;
        rom_memory[26910] = 3'b110;
        rom_memory[26911] = 3'b110;
        rom_memory[26912] = 3'b111;
        rom_memory[26913] = 3'b111;
        rom_memory[26914] = 3'b111;
        rom_memory[26915] = 3'b111;
        rom_memory[26916] = 3'b111;
        rom_memory[26917] = 3'b111;
        rom_memory[26918] = 3'b111;
        rom_memory[26919] = 3'b111;
        rom_memory[26920] = 3'b110;
        rom_memory[26921] = 3'b110;
        rom_memory[26922] = 3'b110;
        rom_memory[26923] = 3'b111;
        rom_memory[26924] = 3'b111;
        rom_memory[26925] = 3'b111;
        rom_memory[26926] = 3'b111;
        rom_memory[26927] = 3'b111;
        rom_memory[26928] = 3'b111;
        rom_memory[26929] = 3'b111;
        rom_memory[26930] = 3'b111;
        rom_memory[26931] = 3'b111;
        rom_memory[26932] = 3'b111;
        rom_memory[26933] = 3'b111;
        rom_memory[26934] = 3'b111;
        rom_memory[26935] = 3'b111;
        rom_memory[26936] = 3'b111;
        rom_memory[26937] = 3'b111;
        rom_memory[26938] = 3'b111;
        rom_memory[26939] = 3'b110;
        rom_memory[26940] = 3'b110;
        rom_memory[26941] = 3'b100;
        rom_memory[26942] = 3'b110;
        rom_memory[26943] = 3'b110;
        rom_memory[26944] = 3'b110;
        rom_memory[26945] = 3'b110;
        rom_memory[26946] = 3'b110;
        rom_memory[26947] = 3'b100;
        rom_memory[26948] = 3'b100;
        rom_memory[26949] = 3'b100;
        rom_memory[26950] = 3'b110;
        rom_memory[26951] = 3'b110;
        rom_memory[26952] = 3'b110;
        rom_memory[26953] = 3'b110;
        rom_memory[26954] = 3'b110;
        rom_memory[26955] = 3'b110;
        rom_memory[26956] = 3'b110;
        rom_memory[26957] = 3'b110;
        rom_memory[26958] = 3'b110;
        rom_memory[26959] = 3'b110;
        rom_memory[26960] = 3'b110;
        rom_memory[26961] = 3'b110;
        rom_memory[26962] = 3'b110;
        rom_memory[26963] = 3'b110;
        rom_memory[26964] = 3'b110;
        rom_memory[26965] = 3'b110;
        rom_memory[26966] = 3'b110;
        rom_memory[26967] = 3'b110;
        rom_memory[26968] = 3'b110;
        rom_memory[26969] = 3'b110;
        rom_memory[26970] = 3'b110;
        rom_memory[26971] = 3'b110;
        rom_memory[26972] = 3'b110;
        rom_memory[26973] = 3'b110;
        rom_memory[26974] = 3'b110;
        rom_memory[26975] = 3'b110;
        rom_memory[26976] = 3'b110;
        rom_memory[26977] = 3'b110;
        rom_memory[26978] = 3'b110;
        rom_memory[26979] = 3'b110;
        rom_memory[26980] = 3'b110;
        rom_memory[26981] = 3'b110;
        rom_memory[26982] = 3'b110;
        rom_memory[26983] = 3'b110;
        rom_memory[26984] = 3'b110;
        rom_memory[26985] = 3'b110;
        rom_memory[26986] = 3'b110;
        rom_memory[26987] = 3'b110;
        rom_memory[26988] = 3'b110;
        rom_memory[26989] = 3'b110;
        rom_memory[26990] = 3'b110;
        rom_memory[26991] = 3'b110;
        rom_memory[26992] = 3'b110;
        rom_memory[26993] = 3'b110;
        rom_memory[26994] = 3'b110;
        rom_memory[26995] = 3'b110;
        rom_memory[26996] = 3'b110;
        rom_memory[26997] = 3'b110;
        rom_memory[26998] = 3'b110;
        rom_memory[26999] = 3'b110;
        rom_memory[27000] = 3'b110;
        rom_memory[27001] = 3'b110;
        rom_memory[27002] = 3'b110;
        rom_memory[27003] = 3'b100;
        rom_memory[27004] = 3'b000;
        rom_memory[27005] = 3'b100;
        rom_memory[27006] = 3'b100;
        rom_memory[27007] = 3'b000;
        rom_memory[27008] = 3'b000;
        rom_memory[27009] = 3'b000;
        rom_memory[27010] = 3'b000;
        rom_memory[27011] = 3'b000;
        rom_memory[27012] = 3'b000;
        rom_memory[27013] = 3'b000;
        rom_memory[27014] = 3'b111;
        rom_memory[27015] = 3'b110;
        rom_memory[27016] = 3'b110;
        rom_memory[27017] = 3'b110;
        rom_memory[27018] = 3'b110;
        rom_memory[27019] = 3'b110;
        rom_memory[27020] = 3'b110;
        rom_memory[27021] = 3'b110;
        rom_memory[27022] = 3'b110;
        rom_memory[27023] = 3'b110;
        rom_memory[27024] = 3'b110;
        rom_memory[27025] = 3'b110;
        rom_memory[27026] = 3'b110;
        rom_memory[27027] = 3'b110;
        rom_memory[27028] = 3'b110;
        rom_memory[27029] = 3'b110;
        rom_memory[27030] = 3'b110;
        rom_memory[27031] = 3'b110;
        rom_memory[27032] = 3'b110;
        rom_memory[27033] = 3'b110;
        rom_memory[27034] = 3'b110;
        rom_memory[27035] = 3'b110;
        rom_memory[27036] = 3'b110;
        rom_memory[27037] = 3'b110;
        rom_memory[27038] = 3'b110;
        rom_memory[27039] = 3'b110;
        rom_memory[27040] = 3'b110;
        rom_memory[27041] = 3'b110;
        rom_memory[27042] = 3'b110;
        rom_memory[27043] = 3'b110;
        rom_memory[27044] = 3'b110;
        rom_memory[27045] = 3'b110;
        rom_memory[27046] = 3'b110;
        rom_memory[27047] = 3'b110;
        rom_memory[27048] = 3'b110;
        rom_memory[27049] = 3'b110;
        rom_memory[27050] = 3'b111;
        rom_memory[27051] = 3'b110;
        rom_memory[27052] = 3'b110;
        rom_memory[27053] = 3'b111;
        rom_memory[27054] = 3'b110;
        rom_memory[27055] = 3'b110;
        rom_memory[27056] = 3'b110;
        rom_memory[27057] = 3'b111;
        rom_memory[27058] = 3'b111;
        rom_memory[27059] = 3'b111;
        rom_memory[27060] = 3'b110;
        rom_memory[27061] = 3'b110;
        rom_memory[27062] = 3'b111;
        rom_memory[27063] = 3'b111;
        rom_memory[27064] = 3'b111;
        rom_memory[27065] = 3'b111;
        rom_memory[27066] = 3'b111;
        rom_memory[27067] = 3'b111;
        rom_memory[27068] = 3'b111;
        rom_memory[27069] = 3'b111;
        rom_memory[27070] = 3'b111;
        rom_memory[27071] = 3'b111;
        rom_memory[27072] = 3'b111;
        rom_memory[27073] = 3'b111;
        rom_memory[27074] = 3'b111;
        rom_memory[27075] = 3'b111;
        rom_memory[27076] = 3'b111;
        rom_memory[27077] = 3'b111;
        rom_memory[27078] = 3'b111;
        rom_memory[27079] = 3'b111;
        rom_memory[27080] = 3'b111;
        rom_memory[27081] = 3'b111;
        rom_memory[27082] = 3'b111;
        rom_memory[27083] = 3'b111;
        rom_memory[27084] = 3'b111;
        rom_memory[27085] = 3'b111;
        rom_memory[27086] = 3'b111;
        rom_memory[27087] = 3'b111;
        rom_memory[27088] = 3'b111;
        rom_memory[27089] = 3'b111;
        rom_memory[27090] = 3'b111;
        rom_memory[27091] = 3'b111;
        rom_memory[27092] = 3'b111;
        rom_memory[27093] = 3'b111;
        rom_memory[27094] = 3'b111;
        rom_memory[27095] = 3'b111;
        rom_memory[27096] = 3'b111;
        rom_memory[27097] = 3'b111;
        rom_memory[27098] = 3'b111;
        rom_memory[27099] = 3'b111;
        rom_memory[27100] = 3'b111;
        rom_memory[27101] = 3'b111;
        rom_memory[27102] = 3'b111;
        rom_memory[27103] = 3'b111;
        rom_memory[27104] = 3'b111;
        rom_memory[27105] = 3'b111;
        rom_memory[27106] = 3'b111;
        rom_memory[27107] = 3'b111;
        rom_memory[27108] = 3'b111;
        rom_memory[27109] = 3'b111;
        rom_memory[27110] = 3'b111;
        rom_memory[27111] = 3'b111;
        rom_memory[27112] = 3'b111;
        rom_memory[27113] = 3'b111;
        rom_memory[27114] = 3'b111;
        rom_memory[27115] = 3'b111;
        rom_memory[27116] = 3'b111;
        rom_memory[27117] = 3'b111;
        rom_memory[27118] = 3'b111;
        rom_memory[27119] = 3'b111;
        rom_memory[27120] = 3'b110;
        rom_memory[27121] = 3'b110;
        rom_memory[27122] = 3'b110;
        rom_memory[27123] = 3'b110;
        rom_memory[27124] = 3'b110;
        rom_memory[27125] = 3'b110;
        rom_memory[27126] = 3'b110;
        rom_memory[27127] = 3'b110;
        rom_memory[27128] = 3'b110;
        rom_memory[27129] = 3'b110;
        rom_memory[27130] = 3'b110;
        rom_memory[27131] = 3'b110;
        rom_memory[27132] = 3'b110;
        rom_memory[27133] = 3'b110;
        rom_memory[27134] = 3'b110;
        rom_memory[27135] = 3'b110;
        rom_memory[27136] = 3'b111;
        rom_memory[27137] = 3'b111;
        rom_memory[27138] = 3'b111;
        rom_memory[27139] = 3'b110;
        rom_memory[27140] = 3'b110;
        rom_memory[27141] = 3'b110;
        rom_memory[27142] = 3'b110;
        rom_memory[27143] = 3'b110;
        rom_memory[27144] = 3'b110;
        rom_memory[27145] = 3'b110;
        rom_memory[27146] = 3'b110;
        rom_memory[27147] = 3'b110;
        rom_memory[27148] = 3'b110;
        rom_memory[27149] = 3'b110;
        rom_memory[27150] = 3'b110;
        rom_memory[27151] = 3'b110;
        rom_memory[27152] = 3'b111;
        rom_memory[27153] = 3'b111;
        rom_memory[27154] = 3'b111;
        rom_memory[27155] = 3'b111;
        rom_memory[27156] = 3'b111;
        rom_memory[27157] = 3'b110;
        rom_memory[27158] = 3'b110;
        rom_memory[27159] = 3'b110;
        rom_memory[27160] = 3'b110;
        rom_memory[27161] = 3'b110;
        rom_memory[27162] = 3'b110;
        rom_memory[27163] = 3'b110;
        rom_memory[27164] = 3'b110;
        rom_memory[27165] = 3'b110;
        rom_memory[27166] = 3'b111;
        rom_memory[27167] = 3'b110;
        rom_memory[27168] = 3'b110;
        rom_memory[27169] = 3'b110;
        rom_memory[27170] = 3'b111;
        rom_memory[27171] = 3'b111;
        rom_memory[27172] = 3'b111;
        rom_memory[27173] = 3'b111;
        rom_memory[27174] = 3'b111;
        rom_memory[27175] = 3'b111;
        rom_memory[27176] = 3'b111;
        rom_memory[27177] = 3'b111;
        rom_memory[27178] = 3'b111;
        rom_memory[27179] = 3'b110;
        rom_memory[27180] = 3'b110;
        rom_memory[27181] = 3'b110;
        rom_memory[27182] = 3'b100;
        rom_memory[27183] = 3'b110;
        rom_memory[27184] = 3'b110;
        rom_memory[27185] = 3'b110;
        rom_memory[27186] = 3'b110;
        rom_memory[27187] = 3'b100;
        rom_memory[27188] = 3'b100;
        rom_memory[27189] = 3'b100;
        rom_memory[27190] = 3'b100;
        rom_memory[27191] = 3'b100;
        rom_memory[27192] = 3'b100;
        rom_memory[27193] = 3'b110;
        rom_memory[27194] = 3'b110;
        rom_memory[27195] = 3'b110;
        rom_memory[27196] = 3'b110;
        rom_memory[27197] = 3'b110;
        rom_memory[27198] = 3'b110;
        rom_memory[27199] = 3'b110;
        rom_memory[27200] = 3'b110;
        rom_memory[27201] = 3'b110;
        rom_memory[27202] = 3'b110;
        rom_memory[27203] = 3'b110;
        rom_memory[27204] = 3'b110;
        rom_memory[27205] = 3'b110;
        rom_memory[27206] = 3'b110;
        rom_memory[27207] = 3'b110;
        rom_memory[27208] = 3'b110;
        rom_memory[27209] = 3'b110;
        rom_memory[27210] = 3'b110;
        rom_memory[27211] = 3'b110;
        rom_memory[27212] = 3'b110;
        rom_memory[27213] = 3'b110;
        rom_memory[27214] = 3'b110;
        rom_memory[27215] = 3'b110;
        rom_memory[27216] = 3'b110;
        rom_memory[27217] = 3'b110;
        rom_memory[27218] = 3'b110;
        rom_memory[27219] = 3'b110;
        rom_memory[27220] = 3'b110;
        rom_memory[27221] = 3'b110;
        rom_memory[27222] = 3'b110;
        rom_memory[27223] = 3'b110;
        rom_memory[27224] = 3'b110;
        rom_memory[27225] = 3'b110;
        rom_memory[27226] = 3'b110;
        rom_memory[27227] = 3'b110;
        rom_memory[27228] = 3'b110;
        rom_memory[27229] = 3'b110;
        rom_memory[27230] = 3'b110;
        rom_memory[27231] = 3'b110;
        rom_memory[27232] = 3'b110;
        rom_memory[27233] = 3'b110;
        rom_memory[27234] = 3'b110;
        rom_memory[27235] = 3'b110;
        rom_memory[27236] = 3'b110;
        rom_memory[27237] = 3'b110;
        rom_memory[27238] = 3'b110;
        rom_memory[27239] = 3'b110;
        rom_memory[27240] = 3'b110;
        rom_memory[27241] = 3'b110;
        rom_memory[27242] = 3'b110;
        rom_memory[27243] = 3'b110;
        rom_memory[27244] = 3'b100;
        rom_memory[27245] = 3'b100;
        rom_memory[27246] = 3'b100;
        rom_memory[27247] = 3'b100;
        rom_memory[27248] = 3'b000;
        rom_memory[27249] = 3'b000;
        rom_memory[27250] = 3'b000;
        rom_memory[27251] = 3'b000;
        rom_memory[27252] = 3'b000;
        rom_memory[27253] = 3'b000;
        rom_memory[27254] = 3'b110;
        rom_memory[27255] = 3'b110;
        rom_memory[27256] = 3'b110;
        rom_memory[27257] = 3'b110;
        rom_memory[27258] = 3'b110;
        rom_memory[27259] = 3'b110;
        rom_memory[27260] = 3'b110;
        rom_memory[27261] = 3'b110;
        rom_memory[27262] = 3'b110;
        rom_memory[27263] = 3'b110;
        rom_memory[27264] = 3'b110;
        rom_memory[27265] = 3'b110;
        rom_memory[27266] = 3'b110;
        rom_memory[27267] = 3'b110;
        rom_memory[27268] = 3'b110;
        rom_memory[27269] = 3'b110;
        rom_memory[27270] = 3'b110;
        rom_memory[27271] = 3'b110;
        rom_memory[27272] = 3'b110;
        rom_memory[27273] = 3'b110;
        rom_memory[27274] = 3'b110;
        rom_memory[27275] = 3'b110;
        rom_memory[27276] = 3'b110;
        rom_memory[27277] = 3'b110;
        rom_memory[27278] = 3'b110;
        rom_memory[27279] = 3'b110;
        rom_memory[27280] = 3'b110;
        rom_memory[27281] = 3'b110;
        rom_memory[27282] = 3'b110;
        rom_memory[27283] = 3'b110;
        rom_memory[27284] = 3'b110;
        rom_memory[27285] = 3'b110;
        rom_memory[27286] = 3'b110;
        rom_memory[27287] = 3'b110;
        rom_memory[27288] = 3'b110;
        rom_memory[27289] = 3'b110;
        rom_memory[27290] = 3'b110;
        rom_memory[27291] = 3'b110;
        rom_memory[27292] = 3'b110;
        rom_memory[27293] = 3'b111;
        rom_memory[27294] = 3'b110;
        rom_memory[27295] = 3'b110;
        rom_memory[27296] = 3'b110;
        rom_memory[27297] = 3'b111;
        rom_memory[27298] = 3'b111;
        rom_memory[27299] = 3'b111;
        rom_memory[27300] = 3'b111;
        rom_memory[27301] = 3'b110;
        rom_memory[27302] = 3'b111;
        rom_memory[27303] = 3'b111;
        rom_memory[27304] = 3'b111;
        rom_memory[27305] = 3'b111;
        rom_memory[27306] = 3'b111;
        rom_memory[27307] = 3'b111;
        rom_memory[27308] = 3'b111;
        rom_memory[27309] = 3'b111;
        rom_memory[27310] = 3'b111;
        rom_memory[27311] = 3'b111;
        rom_memory[27312] = 3'b111;
        rom_memory[27313] = 3'b111;
        rom_memory[27314] = 3'b111;
        rom_memory[27315] = 3'b111;
        rom_memory[27316] = 3'b111;
        rom_memory[27317] = 3'b111;
        rom_memory[27318] = 3'b111;
        rom_memory[27319] = 3'b111;
        rom_memory[27320] = 3'b111;
        rom_memory[27321] = 3'b111;
        rom_memory[27322] = 3'b111;
        rom_memory[27323] = 3'b111;
        rom_memory[27324] = 3'b111;
        rom_memory[27325] = 3'b111;
        rom_memory[27326] = 3'b111;
        rom_memory[27327] = 3'b111;
        rom_memory[27328] = 3'b111;
        rom_memory[27329] = 3'b111;
        rom_memory[27330] = 3'b111;
        rom_memory[27331] = 3'b111;
        rom_memory[27332] = 3'b111;
        rom_memory[27333] = 3'b111;
        rom_memory[27334] = 3'b111;
        rom_memory[27335] = 3'b111;
        rom_memory[27336] = 3'b111;
        rom_memory[27337] = 3'b111;
        rom_memory[27338] = 3'b111;
        rom_memory[27339] = 3'b111;
        rom_memory[27340] = 3'b111;
        rom_memory[27341] = 3'b111;
        rom_memory[27342] = 3'b111;
        rom_memory[27343] = 3'b111;
        rom_memory[27344] = 3'b111;
        rom_memory[27345] = 3'b111;
        rom_memory[27346] = 3'b111;
        rom_memory[27347] = 3'b111;
        rom_memory[27348] = 3'b111;
        rom_memory[27349] = 3'b111;
        rom_memory[27350] = 3'b111;
        rom_memory[27351] = 3'b111;
        rom_memory[27352] = 3'b111;
        rom_memory[27353] = 3'b111;
        rom_memory[27354] = 3'b111;
        rom_memory[27355] = 3'b111;
        rom_memory[27356] = 3'b111;
        rom_memory[27357] = 3'b111;
        rom_memory[27358] = 3'b111;
        rom_memory[27359] = 3'b111;
        rom_memory[27360] = 3'b110;
        rom_memory[27361] = 3'b110;
        rom_memory[27362] = 3'b110;
        rom_memory[27363] = 3'b110;
        rom_memory[27364] = 3'b110;
        rom_memory[27365] = 3'b110;
        rom_memory[27366] = 3'b110;
        rom_memory[27367] = 3'b110;
        rom_memory[27368] = 3'b110;
        rom_memory[27369] = 3'b110;
        rom_memory[27370] = 3'b110;
        rom_memory[27371] = 3'b110;
        rom_memory[27372] = 3'b110;
        rom_memory[27373] = 3'b110;
        rom_memory[27374] = 3'b110;
        rom_memory[27375] = 3'b111;
        rom_memory[27376] = 3'b111;
        rom_memory[27377] = 3'b111;
        rom_memory[27378] = 3'b111;
        rom_memory[27379] = 3'b111;
        rom_memory[27380] = 3'b111;
        rom_memory[27381] = 3'b110;
        rom_memory[27382] = 3'b111;
        rom_memory[27383] = 3'b110;
        rom_memory[27384] = 3'b110;
        rom_memory[27385] = 3'b110;
        rom_memory[27386] = 3'b110;
        rom_memory[27387] = 3'b110;
        rom_memory[27388] = 3'b110;
        rom_memory[27389] = 3'b110;
        rom_memory[27390] = 3'b110;
        rom_memory[27391] = 3'b110;
        rom_memory[27392] = 3'b110;
        rom_memory[27393] = 3'b110;
        rom_memory[27394] = 3'b111;
        rom_memory[27395] = 3'b111;
        rom_memory[27396] = 3'b110;
        rom_memory[27397] = 3'b110;
        rom_memory[27398] = 3'b110;
        rom_memory[27399] = 3'b110;
        rom_memory[27400] = 3'b110;
        rom_memory[27401] = 3'b110;
        rom_memory[27402] = 3'b110;
        rom_memory[27403] = 3'b110;
        rom_memory[27404] = 3'b110;
        rom_memory[27405] = 3'b110;
        rom_memory[27406] = 3'b110;
        rom_memory[27407] = 3'b110;
        rom_memory[27408] = 3'b110;
        rom_memory[27409] = 3'b110;
        rom_memory[27410] = 3'b110;
        rom_memory[27411] = 3'b111;
        rom_memory[27412] = 3'b111;
        rom_memory[27413] = 3'b111;
        rom_memory[27414] = 3'b111;
        rom_memory[27415] = 3'b111;
        rom_memory[27416] = 3'b111;
        rom_memory[27417] = 3'b111;
        rom_memory[27418] = 3'b111;
        rom_memory[27419] = 3'b111;
        rom_memory[27420] = 3'b110;
        rom_memory[27421] = 3'b110;
        rom_memory[27422] = 3'b110;
        rom_memory[27423] = 3'b100;
        rom_memory[27424] = 3'b110;
        rom_memory[27425] = 3'b110;
        rom_memory[27426] = 3'b100;
        rom_memory[27427] = 3'b100;
        rom_memory[27428] = 3'b100;
        rom_memory[27429] = 3'b100;
        rom_memory[27430] = 3'b100;
        rom_memory[27431] = 3'b100;
        rom_memory[27432] = 3'b100;
        rom_memory[27433] = 3'b110;
        rom_memory[27434] = 3'b110;
        rom_memory[27435] = 3'b110;
        rom_memory[27436] = 3'b110;
        rom_memory[27437] = 3'b110;
        rom_memory[27438] = 3'b110;
        rom_memory[27439] = 3'b110;
        rom_memory[27440] = 3'b110;
        rom_memory[27441] = 3'b110;
        rom_memory[27442] = 3'b110;
        rom_memory[27443] = 3'b110;
        rom_memory[27444] = 3'b110;
        rom_memory[27445] = 3'b110;
        rom_memory[27446] = 3'b110;
        rom_memory[27447] = 3'b110;
        rom_memory[27448] = 3'b110;
        rom_memory[27449] = 3'b110;
        rom_memory[27450] = 3'b110;
        rom_memory[27451] = 3'b110;
        rom_memory[27452] = 3'b110;
        rom_memory[27453] = 3'b110;
        rom_memory[27454] = 3'b110;
        rom_memory[27455] = 3'b110;
        rom_memory[27456] = 3'b110;
        rom_memory[27457] = 3'b110;
        rom_memory[27458] = 3'b110;
        rom_memory[27459] = 3'b110;
        rom_memory[27460] = 3'b110;
        rom_memory[27461] = 3'b110;
        rom_memory[27462] = 3'b110;
        rom_memory[27463] = 3'b110;
        rom_memory[27464] = 3'b110;
        rom_memory[27465] = 3'b110;
        rom_memory[27466] = 3'b110;
        rom_memory[27467] = 3'b110;
        rom_memory[27468] = 3'b110;
        rom_memory[27469] = 3'b110;
        rom_memory[27470] = 3'b110;
        rom_memory[27471] = 3'b110;
        rom_memory[27472] = 3'b110;
        rom_memory[27473] = 3'b110;
        rom_memory[27474] = 3'b110;
        rom_memory[27475] = 3'b110;
        rom_memory[27476] = 3'b110;
        rom_memory[27477] = 3'b110;
        rom_memory[27478] = 3'b110;
        rom_memory[27479] = 3'b110;
        rom_memory[27480] = 3'b110;
        rom_memory[27481] = 3'b110;
        rom_memory[27482] = 3'b110;
        rom_memory[27483] = 3'b110;
        rom_memory[27484] = 3'b110;
        rom_memory[27485] = 3'b110;
        rom_memory[27486] = 3'b100;
        rom_memory[27487] = 3'b110;
        rom_memory[27488] = 3'b100;
        rom_memory[27489] = 3'b000;
        rom_memory[27490] = 3'b000;
        rom_memory[27491] = 3'b000;
        rom_memory[27492] = 3'b000;
        rom_memory[27493] = 3'b000;
        rom_memory[27494] = 3'b100;
        rom_memory[27495] = 3'b110;
        rom_memory[27496] = 3'b110;
        rom_memory[27497] = 3'b110;
        rom_memory[27498] = 3'b110;
        rom_memory[27499] = 3'b110;
        rom_memory[27500] = 3'b110;
        rom_memory[27501] = 3'b110;
        rom_memory[27502] = 3'b110;
        rom_memory[27503] = 3'b110;
        rom_memory[27504] = 3'b110;
        rom_memory[27505] = 3'b110;
        rom_memory[27506] = 3'b110;
        rom_memory[27507] = 3'b110;
        rom_memory[27508] = 3'b110;
        rom_memory[27509] = 3'b110;
        rom_memory[27510] = 3'b110;
        rom_memory[27511] = 3'b110;
        rom_memory[27512] = 3'b110;
        rom_memory[27513] = 3'b110;
        rom_memory[27514] = 3'b110;
        rom_memory[27515] = 3'b110;
        rom_memory[27516] = 3'b110;
        rom_memory[27517] = 3'b110;
        rom_memory[27518] = 3'b110;
        rom_memory[27519] = 3'b110;
        rom_memory[27520] = 3'b110;
        rom_memory[27521] = 3'b110;
        rom_memory[27522] = 3'b110;
        rom_memory[27523] = 3'b110;
        rom_memory[27524] = 3'b110;
        rom_memory[27525] = 3'b110;
        rom_memory[27526] = 3'b110;
        rom_memory[27527] = 3'b110;
        rom_memory[27528] = 3'b110;
        rom_memory[27529] = 3'b110;
        rom_memory[27530] = 3'b110;
        rom_memory[27531] = 3'b110;
        rom_memory[27532] = 3'b110;
        rom_memory[27533] = 3'b110;
        rom_memory[27534] = 3'b110;
        rom_memory[27535] = 3'b110;
        rom_memory[27536] = 3'b110;
        rom_memory[27537] = 3'b111;
        rom_memory[27538] = 3'b111;
        rom_memory[27539] = 3'b111;
        rom_memory[27540] = 3'b111;
        rom_memory[27541] = 3'b110;
        rom_memory[27542] = 3'b111;
        rom_memory[27543] = 3'b111;
        rom_memory[27544] = 3'b111;
        rom_memory[27545] = 3'b111;
        rom_memory[27546] = 3'b111;
        rom_memory[27547] = 3'b111;
        rom_memory[27548] = 3'b111;
        rom_memory[27549] = 3'b111;
        rom_memory[27550] = 3'b111;
        rom_memory[27551] = 3'b111;
        rom_memory[27552] = 3'b111;
        rom_memory[27553] = 3'b111;
        rom_memory[27554] = 3'b111;
        rom_memory[27555] = 3'b111;
        rom_memory[27556] = 3'b111;
        rom_memory[27557] = 3'b111;
        rom_memory[27558] = 3'b111;
        rom_memory[27559] = 3'b111;
        rom_memory[27560] = 3'b111;
        rom_memory[27561] = 3'b111;
        rom_memory[27562] = 3'b111;
        rom_memory[27563] = 3'b111;
        rom_memory[27564] = 3'b111;
        rom_memory[27565] = 3'b111;
        rom_memory[27566] = 3'b111;
        rom_memory[27567] = 3'b111;
        rom_memory[27568] = 3'b111;
        rom_memory[27569] = 3'b111;
        rom_memory[27570] = 3'b111;
        rom_memory[27571] = 3'b111;
        rom_memory[27572] = 3'b111;
        rom_memory[27573] = 3'b111;
        rom_memory[27574] = 3'b111;
        rom_memory[27575] = 3'b111;
        rom_memory[27576] = 3'b111;
        rom_memory[27577] = 3'b111;
        rom_memory[27578] = 3'b111;
        rom_memory[27579] = 3'b111;
        rom_memory[27580] = 3'b111;
        rom_memory[27581] = 3'b111;
        rom_memory[27582] = 3'b111;
        rom_memory[27583] = 3'b111;
        rom_memory[27584] = 3'b111;
        rom_memory[27585] = 3'b111;
        rom_memory[27586] = 3'b111;
        rom_memory[27587] = 3'b111;
        rom_memory[27588] = 3'b111;
        rom_memory[27589] = 3'b111;
        rom_memory[27590] = 3'b111;
        rom_memory[27591] = 3'b111;
        rom_memory[27592] = 3'b111;
        rom_memory[27593] = 3'b111;
        rom_memory[27594] = 3'b111;
        rom_memory[27595] = 3'b111;
        rom_memory[27596] = 3'b111;
        rom_memory[27597] = 3'b111;
        rom_memory[27598] = 3'b111;
        rom_memory[27599] = 3'b111;
        rom_memory[27600] = 3'b110;
        rom_memory[27601] = 3'b110;
        rom_memory[27602] = 3'b110;
        rom_memory[27603] = 3'b110;
        rom_memory[27604] = 3'b110;
        rom_memory[27605] = 3'b110;
        rom_memory[27606] = 3'b110;
        rom_memory[27607] = 3'b110;
        rom_memory[27608] = 3'b110;
        rom_memory[27609] = 3'b110;
        rom_memory[27610] = 3'b110;
        rom_memory[27611] = 3'b110;
        rom_memory[27612] = 3'b110;
        rom_memory[27613] = 3'b111;
        rom_memory[27614] = 3'b111;
        rom_memory[27615] = 3'b111;
        rom_memory[27616] = 3'b111;
        rom_memory[27617] = 3'b111;
        rom_memory[27618] = 3'b111;
        rom_memory[27619] = 3'b111;
        rom_memory[27620] = 3'b111;
        rom_memory[27621] = 3'b111;
        rom_memory[27622] = 3'b111;
        rom_memory[27623] = 3'b111;
        rom_memory[27624] = 3'b110;
        rom_memory[27625] = 3'b110;
        rom_memory[27626] = 3'b110;
        rom_memory[27627] = 3'b110;
        rom_memory[27628] = 3'b110;
        rom_memory[27629] = 3'b110;
        rom_memory[27630] = 3'b110;
        rom_memory[27631] = 3'b110;
        rom_memory[27632] = 3'b110;
        rom_memory[27633] = 3'b110;
        rom_memory[27634] = 3'b111;
        rom_memory[27635] = 3'b111;
        rom_memory[27636] = 3'b111;
        rom_memory[27637] = 3'b110;
        rom_memory[27638] = 3'b110;
        rom_memory[27639] = 3'b110;
        rom_memory[27640] = 3'b110;
        rom_memory[27641] = 3'b110;
        rom_memory[27642] = 3'b110;
        rom_memory[27643] = 3'b110;
        rom_memory[27644] = 3'b110;
        rom_memory[27645] = 3'b110;
        rom_memory[27646] = 3'b110;
        rom_memory[27647] = 3'b110;
        rom_memory[27648] = 3'b110;
        rom_memory[27649] = 3'b110;
        rom_memory[27650] = 3'b110;
        rom_memory[27651] = 3'b110;
        rom_memory[27652] = 3'b111;
        rom_memory[27653] = 3'b111;
        rom_memory[27654] = 3'b111;
        rom_memory[27655] = 3'b111;
        rom_memory[27656] = 3'b111;
        rom_memory[27657] = 3'b111;
        rom_memory[27658] = 3'b111;
        rom_memory[27659] = 3'b111;
        rom_memory[27660] = 3'b111;
        rom_memory[27661] = 3'b110;
        rom_memory[27662] = 3'b110;
        rom_memory[27663] = 3'b100;
        rom_memory[27664] = 3'b110;
        rom_memory[27665] = 3'b110;
        rom_memory[27666] = 3'b100;
        rom_memory[27667] = 3'b100;
        rom_memory[27668] = 3'b100;
        rom_memory[27669] = 3'b100;
        rom_memory[27670] = 3'b100;
        rom_memory[27671] = 3'b100;
        rom_memory[27672] = 3'b100;
        rom_memory[27673] = 3'b100;
        rom_memory[27674] = 3'b110;
        rom_memory[27675] = 3'b110;
        rom_memory[27676] = 3'b110;
        rom_memory[27677] = 3'b110;
        rom_memory[27678] = 3'b110;
        rom_memory[27679] = 3'b110;
        rom_memory[27680] = 3'b110;
        rom_memory[27681] = 3'b110;
        rom_memory[27682] = 3'b110;
        rom_memory[27683] = 3'b110;
        rom_memory[27684] = 3'b110;
        rom_memory[27685] = 3'b110;
        rom_memory[27686] = 3'b110;
        rom_memory[27687] = 3'b110;
        rom_memory[27688] = 3'b110;
        rom_memory[27689] = 3'b110;
        rom_memory[27690] = 3'b110;
        rom_memory[27691] = 3'b110;
        rom_memory[27692] = 3'b110;
        rom_memory[27693] = 3'b110;
        rom_memory[27694] = 3'b110;
        rom_memory[27695] = 3'b110;
        rom_memory[27696] = 3'b110;
        rom_memory[27697] = 3'b110;
        rom_memory[27698] = 3'b100;
        rom_memory[27699] = 3'b110;
        rom_memory[27700] = 3'b110;
        rom_memory[27701] = 3'b110;
        rom_memory[27702] = 3'b110;
        rom_memory[27703] = 3'b110;
        rom_memory[27704] = 3'b110;
        rom_memory[27705] = 3'b110;
        rom_memory[27706] = 3'b110;
        rom_memory[27707] = 3'b110;
        rom_memory[27708] = 3'b110;
        rom_memory[27709] = 3'b110;
        rom_memory[27710] = 3'b110;
        rom_memory[27711] = 3'b110;
        rom_memory[27712] = 3'b110;
        rom_memory[27713] = 3'b110;
        rom_memory[27714] = 3'b110;
        rom_memory[27715] = 3'b110;
        rom_memory[27716] = 3'b110;
        rom_memory[27717] = 3'b110;
        rom_memory[27718] = 3'b110;
        rom_memory[27719] = 3'b110;
        rom_memory[27720] = 3'b110;
        rom_memory[27721] = 3'b110;
        rom_memory[27722] = 3'b100;
        rom_memory[27723] = 3'b110;
        rom_memory[27724] = 3'b110;
        rom_memory[27725] = 3'b110;
        rom_memory[27726] = 3'b110;
        rom_memory[27727] = 3'b110;
        rom_memory[27728] = 3'b110;
        rom_memory[27729] = 3'b000;
        rom_memory[27730] = 3'b000;
        rom_memory[27731] = 3'b000;
        rom_memory[27732] = 3'b000;
        rom_memory[27733] = 3'b000;
        rom_memory[27734] = 3'b000;
        rom_memory[27735] = 3'b110;
        rom_memory[27736] = 3'b110;
        rom_memory[27737] = 3'b110;
        rom_memory[27738] = 3'b110;
        rom_memory[27739] = 3'b110;
        rom_memory[27740] = 3'b110;
        rom_memory[27741] = 3'b110;
        rom_memory[27742] = 3'b110;
        rom_memory[27743] = 3'b110;
        rom_memory[27744] = 3'b110;
        rom_memory[27745] = 3'b110;
        rom_memory[27746] = 3'b110;
        rom_memory[27747] = 3'b110;
        rom_memory[27748] = 3'b110;
        rom_memory[27749] = 3'b110;
        rom_memory[27750] = 3'b110;
        rom_memory[27751] = 3'b110;
        rom_memory[27752] = 3'b110;
        rom_memory[27753] = 3'b110;
        rom_memory[27754] = 3'b110;
        rom_memory[27755] = 3'b110;
        rom_memory[27756] = 3'b110;
        rom_memory[27757] = 3'b110;
        rom_memory[27758] = 3'b110;
        rom_memory[27759] = 3'b110;
        rom_memory[27760] = 3'b110;
        rom_memory[27761] = 3'b110;
        rom_memory[27762] = 3'b110;
        rom_memory[27763] = 3'b110;
        rom_memory[27764] = 3'b110;
        rom_memory[27765] = 3'b110;
        rom_memory[27766] = 3'b110;
        rom_memory[27767] = 3'b110;
        rom_memory[27768] = 3'b110;
        rom_memory[27769] = 3'b110;
        rom_memory[27770] = 3'b110;
        rom_memory[27771] = 3'b110;
        rom_memory[27772] = 3'b111;
        rom_memory[27773] = 3'b110;
        rom_memory[27774] = 3'b110;
        rom_memory[27775] = 3'b110;
        rom_memory[27776] = 3'b110;
        rom_memory[27777] = 3'b111;
        rom_memory[27778] = 3'b111;
        rom_memory[27779] = 3'b110;
        rom_memory[27780] = 3'b110;
        rom_memory[27781] = 3'b111;
        rom_memory[27782] = 3'b111;
        rom_memory[27783] = 3'b111;
        rom_memory[27784] = 3'b111;
        rom_memory[27785] = 3'b111;
        rom_memory[27786] = 3'b111;
        rom_memory[27787] = 3'b111;
        rom_memory[27788] = 3'b111;
        rom_memory[27789] = 3'b111;
        rom_memory[27790] = 3'b111;
        rom_memory[27791] = 3'b111;
        rom_memory[27792] = 3'b111;
        rom_memory[27793] = 3'b111;
        rom_memory[27794] = 3'b111;
        rom_memory[27795] = 3'b111;
        rom_memory[27796] = 3'b111;
        rom_memory[27797] = 3'b111;
        rom_memory[27798] = 3'b111;
        rom_memory[27799] = 3'b111;
        rom_memory[27800] = 3'b111;
        rom_memory[27801] = 3'b111;
        rom_memory[27802] = 3'b111;
        rom_memory[27803] = 3'b111;
        rom_memory[27804] = 3'b111;
        rom_memory[27805] = 3'b111;
        rom_memory[27806] = 3'b111;
        rom_memory[27807] = 3'b111;
        rom_memory[27808] = 3'b111;
        rom_memory[27809] = 3'b111;
        rom_memory[27810] = 3'b111;
        rom_memory[27811] = 3'b111;
        rom_memory[27812] = 3'b111;
        rom_memory[27813] = 3'b111;
        rom_memory[27814] = 3'b111;
        rom_memory[27815] = 3'b111;
        rom_memory[27816] = 3'b111;
        rom_memory[27817] = 3'b111;
        rom_memory[27818] = 3'b111;
        rom_memory[27819] = 3'b111;
        rom_memory[27820] = 3'b111;
        rom_memory[27821] = 3'b111;
        rom_memory[27822] = 3'b111;
        rom_memory[27823] = 3'b111;
        rom_memory[27824] = 3'b111;
        rom_memory[27825] = 3'b111;
        rom_memory[27826] = 3'b111;
        rom_memory[27827] = 3'b111;
        rom_memory[27828] = 3'b111;
        rom_memory[27829] = 3'b111;
        rom_memory[27830] = 3'b111;
        rom_memory[27831] = 3'b111;
        rom_memory[27832] = 3'b111;
        rom_memory[27833] = 3'b111;
        rom_memory[27834] = 3'b111;
        rom_memory[27835] = 3'b111;
        rom_memory[27836] = 3'b111;
        rom_memory[27837] = 3'b111;
        rom_memory[27838] = 3'b111;
        rom_memory[27839] = 3'b111;
        rom_memory[27840] = 3'b110;
        rom_memory[27841] = 3'b110;
        rom_memory[27842] = 3'b110;
        rom_memory[27843] = 3'b110;
        rom_memory[27844] = 3'b110;
        rom_memory[27845] = 3'b110;
        rom_memory[27846] = 3'b110;
        rom_memory[27847] = 3'b110;
        rom_memory[27848] = 3'b110;
        rom_memory[27849] = 3'b110;
        rom_memory[27850] = 3'b110;
        rom_memory[27851] = 3'b110;
        rom_memory[27852] = 3'b111;
        rom_memory[27853] = 3'b111;
        rom_memory[27854] = 3'b111;
        rom_memory[27855] = 3'b111;
        rom_memory[27856] = 3'b111;
        rom_memory[27857] = 3'b111;
        rom_memory[27858] = 3'b111;
        rom_memory[27859] = 3'b111;
        rom_memory[27860] = 3'b111;
        rom_memory[27861] = 3'b111;
        rom_memory[27862] = 3'b111;
        rom_memory[27863] = 3'b111;
        rom_memory[27864] = 3'b111;
        rom_memory[27865] = 3'b111;
        rom_memory[27866] = 3'b110;
        rom_memory[27867] = 3'b110;
        rom_memory[27868] = 3'b110;
        rom_memory[27869] = 3'b110;
        rom_memory[27870] = 3'b110;
        rom_memory[27871] = 3'b110;
        rom_memory[27872] = 3'b110;
        rom_memory[27873] = 3'b110;
        rom_memory[27874] = 3'b111;
        rom_memory[27875] = 3'b111;
        rom_memory[27876] = 3'b110;
        rom_memory[27877] = 3'b110;
        rom_memory[27878] = 3'b110;
        rom_memory[27879] = 3'b110;
        rom_memory[27880] = 3'b110;
        rom_memory[27881] = 3'b110;
        rom_memory[27882] = 3'b110;
        rom_memory[27883] = 3'b110;
        rom_memory[27884] = 3'b110;
        rom_memory[27885] = 3'b110;
        rom_memory[27886] = 3'b110;
        rom_memory[27887] = 3'b110;
        rom_memory[27888] = 3'b110;
        rom_memory[27889] = 3'b110;
        rom_memory[27890] = 3'b110;
        rom_memory[27891] = 3'b110;
        rom_memory[27892] = 3'b111;
        rom_memory[27893] = 3'b111;
        rom_memory[27894] = 3'b111;
        rom_memory[27895] = 3'b111;
        rom_memory[27896] = 3'b111;
        rom_memory[27897] = 3'b111;
        rom_memory[27898] = 3'b111;
        rom_memory[27899] = 3'b111;
        rom_memory[27900] = 3'b111;
        rom_memory[27901] = 3'b111;
        rom_memory[27902] = 3'b110;
        rom_memory[27903] = 3'b110;
        rom_memory[27904] = 3'b100;
        rom_memory[27905] = 3'b110;
        rom_memory[27906] = 3'b110;
        rom_memory[27907] = 3'b100;
        rom_memory[27908] = 3'b100;
        rom_memory[27909] = 3'b100;
        rom_memory[27910] = 3'b100;
        rom_memory[27911] = 3'b100;
        rom_memory[27912] = 3'b100;
        rom_memory[27913] = 3'b100;
        rom_memory[27914] = 3'b100;
        rom_memory[27915] = 3'b110;
        rom_memory[27916] = 3'b110;
        rom_memory[27917] = 3'b110;
        rom_memory[27918] = 3'b110;
        rom_memory[27919] = 3'b110;
        rom_memory[27920] = 3'b110;
        rom_memory[27921] = 3'b110;
        rom_memory[27922] = 3'b110;
        rom_memory[27923] = 3'b110;
        rom_memory[27924] = 3'b110;
        rom_memory[27925] = 3'b110;
        rom_memory[27926] = 3'b110;
        rom_memory[27927] = 3'b110;
        rom_memory[27928] = 3'b110;
        rom_memory[27929] = 3'b110;
        rom_memory[27930] = 3'b110;
        rom_memory[27931] = 3'b110;
        rom_memory[27932] = 3'b110;
        rom_memory[27933] = 3'b110;
        rom_memory[27934] = 3'b110;
        rom_memory[27935] = 3'b110;
        rom_memory[27936] = 3'b110;
        rom_memory[27937] = 3'b110;
        rom_memory[27938] = 3'b100;
        rom_memory[27939] = 3'b110;
        rom_memory[27940] = 3'b110;
        rom_memory[27941] = 3'b110;
        rom_memory[27942] = 3'b110;
        rom_memory[27943] = 3'b110;
        rom_memory[27944] = 3'b110;
        rom_memory[27945] = 3'b110;
        rom_memory[27946] = 3'b110;
        rom_memory[27947] = 3'b110;
        rom_memory[27948] = 3'b110;
        rom_memory[27949] = 3'b110;
        rom_memory[27950] = 3'b110;
        rom_memory[27951] = 3'b110;
        rom_memory[27952] = 3'b110;
        rom_memory[27953] = 3'b110;
        rom_memory[27954] = 3'b110;
        rom_memory[27955] = 3'b110;
        rom_memory[27956] = 3'b110;
        rom_memory[27957] = 3'b110;
        rom_memory[27958] = 3'b110;
        rom_memory[27959] = 3'b110;
        rom_memory[27960] = 3'b110;
        rom_memory[27961] = 3'b110;
        rom_memory[27962] = 3'b100;
        rom_memory[27963] = 3'b110;
        rom_memory[27964] = 3'b110;
        rom_memory[27965] = 3'b110;
        rom_memory[27966] = 3'b110;
        rom_memory[27967] = 3'b110;
        rom_memory[27968] = 3'b110;
        rom_memory[27969] = 3'b110;
        rom_memory[27970] = 3'b000;
        rom_memory[27971] = 3'b000;
        rom_memory[27972] = 3'b000;
        rom_memory[27973] = 3'b000;
        rom_memory[27974] = 3'b000;
        rom_memory[27975] = 3'b100;
        rom_memory[27976] = 3'b110;
        rom_memory[27977] = 3'b110;
        rom_memory[27978] = 3'b110;
        rom_memory[27979] = 3'b110;
        rom_memory[27980] = 3'b110;
        rom_memory[27981] = 3'b110;
        rom_memory[27982] = 3'b110;
        rom_memory[27983] = 3'b110;
        rom_memory[27984] = 3'b110;
        rom_memory[27985] = 3'b110;
        rom_memory[27986] = 3'b110;
        rom_memory[27987] = 3'b110;
        rom_memory[27988] = 3'b110;
        rom_memory[27989] = 3'b110;
        rom_memory[27990] = 3'b110;
        rom_memory[27991] = 3'b110;
        rom_memory[27992] = 3'b110;
        rom_memory[27993] = 3'b110;
        rom_memory[27994] = 3'b110;
        rom_memory[27995] = 3'b110;
        rom_memory[27996] = 3'b110;
        rom_memory[27997] = 3'b110;
        rom_memory[27998] = 3'b110;
        rom_memory[27999] = 3'b110;
        rom_memory[28000] = 3'b110;
        rom_memory[28001] = 3'b110;
        rom_memory[28002] = 3'b110;
        rom_memory[28003] = 3'b110;
        rom_memory[28004] = 3'b110;
        rom_memory[28005] = 3'b110;
        rom_memory[28006] = 3'b110;
        rom_memory[28007] = 3'b110;
        rom_memory[28008] = 3'b110;
        rom_memory[28009] = 3'b110;
        rom_memory[28010] = 3'b110;
        rom_memory[28011] = 3'b110;
        rom_memory[28012] = 3'b110;
        rom_memory[28013] = 3'b110;
        rom_memory[28014] = 3'b110;
        rom_memory[28015] = 3'b110;
        rom_memory[28016] = 3'b110;
        rom_memory[28017] = 3'b110;
        rom_memory[28018] = 3'b111;
        rom_memory[28019] = 3'b110;
        rom_memory[28020] = 3'b110;
        rom_memory[28021] = 3'b110;
        rom_memory[28022] = 3'b110;
        rom_memory[28023] = 3'b111;
        rom_memory[28024] = 3'b111;
        rom_memory[28025] = 3'b111;
        rom_memory[28026] = 3'b111;
        rom_memory[28027] = 3'b111;
        rom_memory[28028] = 3'b111;
        rom_memory[28029] = 3'b111;
        rom_memory[28030] = 3'b111;
        rom_memory[28031] = 3'b111;
        rom_memory[28032] = 3'b111;
        rom_memory[28033] = 3'b111;
        rom_memory[28034] = 3'b111;
        rom_memory[28035] = 3'b111;
        rom_memory[28036] = 3'b111;
        rom_memory[28037] = 3'b111;
        rom_memory[28038] = 3'b111;
        rom_memory[28039] = 3'b111;
        rom_memory[28040] = 3'b111;
        rom_memory[28041] = 3'b111;
        rom_memory[28042] = 3'b111;
        rom_memory[28043] = 3'b111;
        rom_memory[28044] = 3'b111;
        rom_memory[28045] = 3'b111;
        rom_memory[28046] = 3'b111;
        rom_memory[28047] = 3'b111;
        rom_memory[28048] = 3'b111;
        rom_memory[28049] = 3'b111;
        rom_memory[28050] = 3'b111;
        rom_memory[28051] = 3'b111;
        rom_memory[28052] = 3'b111;
        rom_memory[28053] = 3'b111;
        rom_memory[28054] = 3'b111;
        rom_memory[28055] = 3'b111;
        rom_memory[28056] = 3'b111;
        rom_memory[28057] = 3'b111;
        rom_memory[28058] = 3'b111;
        rom_memory[28059] = 3'b111;
        rom_memory[28060] = 3'b111;
        rom_memory[28061] = 3'b111;
        rom_memory[28062] = 3'b111;
        rom_memory[28063] = 3'b111;
        rom_memory[28064] = 3'b111;
        rom_memory[28065] = 3'b111;
        rom_memory[28066] = 3'b111;
        rom_memory[28067] = 3'b111;
        rom_memory[28068] = 3'b111;
        rom_memory[28069] = 3'b111;
        rom_memory[28070] = 3'b111;
        rom_memory[28071] = 3'b111;
        rom_memory[28072] = 3'b111;
        rom_memory[28073] = 3'b111;
        rom_memory[28074] = 3'b111;
        rom_memory[28075] = 3'b111;
        rom_memory[28076] = 3'b111;
        rom_memory[28077] = 3'b111;
        rom_memory[28078] = 3'b111;
        rom_memory[28079] = 3'b111;
        rom_memory[28080] = 3'b110;
        rom_memory[28081] = 3'b110;
        rom_memory[28082] = 3'b110;
        rom_memory[28083] = 3'b110;
        rom_memory[28084] = 3'b110;
        rom_memory[28085] = 3'b110;
        rom_memory[28086] = 3'b110;
        rom_memory[28087] = 3'b110;
        rom_memory[28088] = 3'b110;
        rom_memory[28089] = 3'b110;
        rom_memory[28090] = 3'b110;
        rom_memory[28091] = 3'b110;
        rom_memory[28092] = 3'b111;
        rom_memory[28093] = 3'b111;
        rom_memory[28094] = 3'b111;
        rom_memory[28095] = 3'b111;
        rom_memory[28096] = 3'b111;
        rom_memory[28097] = 3'b111;
        rom_memory[28098] = 3'b111;
        rom_memory[28099] = 3'b111;
        rom_memory[28100] = 3'b111;
        rom_memory[28101] = 3'b111;
        rom_memory[28102] = 3'b111;
        rom_memory[28103] = 3'b111;
        rom_memory[28104] = 3'b111;
        rom_memory[28105] = 3'b111;
        rom_memory[28106] = 3'b110;
        rom_memory[28107] = 3'b110;
        rom_memory[28108] = 3'b110;
        rom_memory[28109] = 3'b110;
        rom_memory[28110] = 3'b110;
        rom_memory[28111] = 3'b110;
        rom_memory[28112] = 3'b110;
        rom_memory[28113] = 3'b110;
        rom_memory[28114] = 3'b111;
        rom_memory[28115] = 3'b111;
        rom_memory[28116] = 3'b110;
        rom_memory[28117] = 3'b110;
        rom_memory[28118] = 3'b110;
        rom_memory[28119] = 3'b110;
        rom_memory[28120] = 3'b110;
        rom_memory[28121] = 3'b110;
        rom_memory[28122] = 3'b110;
        rom_memory[28123] = 3'b110;
        rom_memory[28124] = 3'b110;
        rom_memory[28125] = 3'b110;
        rom_memory[28126] = 3'b110;
        rom_memory[28127] = 3'b110;
        rom_memory[28128] = 3'b110;
        rom_memory[28129] = 3'b110;
        rom_memory[28130] = 3'b110;
        rom_memory[28131] = 3'b110;
        rom_memory[28132] = 3'b111;
        rom_memory[28133] = 3'b111;
        rom_memory[28134] = 3'b111;
        rom_memory[28135] = 3'b111;
        rom_memory[28136] = 3'b111;
        rom_memory[28137] = 3'b111;
        rom_memory[28138] = 3'b111;
        rom_memory[28139] = 3'b111;
        rom_memory[28140] = 3'b111;
        rom_memory[28141] = 3'b111;
        rom_memory[28142] = 3'b111;
        rom_memory[28143] = 3'b110;
        rom_memory[28144] = 3'b110;
        rom_memory[28145] = 3'b100;
        rom_memory[28146] = 3'b110;
        rom_memory[28147] = 3'b110;
        rom_memory[28148] = 3'b100;
        rom_memory[28149] = 3'b100;
        rom_memory[28150] = 3'b100;
        rom_memory[28151] = 3'b100;
        rom_memory[28152] = 3'b100;
        rom_memory[28153] = 3'b100;
        rom_memory[28154] = 3'b100;
        rom_memory[28155] = 3'b100;
        rom_memory[28156] = 3'b110;
        rom_memory[28157] = 3'b110;
        rom_memory[28158] = 3'b110;
        rom_memory[28159] = 3'b110;
        rom_memory[28160] = 3'b110;
        rom_memory[28161] = 3'b110;
        rom_memory[28162] = 3'b110;
        rom_memory[28163] = 3'b110;
        rom_memory[28164] = 3'b110;
        rom_memory[28165] = 3'b110;
        rom_memory[28166] = 3'b110;
        rom_memory[28167] = 3'b110;
        rom_memory[28168] = 3'b110;
        rom_memory[28169] = 3'b110;
        rom_memory[28170] = 3'b110;
        rom_memory[28171] = 3'b110;
        rom_memory[28172] = 3'b110;
        rom_memory[28173] = 3'b110;
        rom_memory[28174] = 3'b110;
        rom_memory[28175] = 3'b110;
        rom_memory[28176] = 3'b110;
        rom_memory[28177] = 3'b110;
        rom_memory[28178] = 3'b110;
        rom_memory[28179] = 3'b110;
        rom_memory[28180] = 3'b110;
        rom_memory[28181] = 3'b110;
        rom_memory[28182] = 3'b110;
        rom_memory[28183] = 3'b110;
        rom_memory[28184] = 3'b110;
        rom_memory[28185] = 3'b110;
        rom_memory[28186] = 3'b110;
        rom_memory[28187] = 3'b110;
        rom_memory[28188] = 3'b110;
        rom_memory[28189] = 3'b110;
        rom_memory[28190] = 3'b110;
        rom_memory[28191] = 3'b110;
        rom_memory[28192] = 3'b110;
        rom_memory[28193] = 3'b110;
        rom_memory[28194] = 3'b110;
        rom_memory[28195] = 3'b110;
        rom_memory[28196] = 3'b110;
        rom_memory[28197] = 3'b110;
        rom_memory[28198] = 3'b110;
        rom_memory[28199] = 3'b110;
        rom_memory[28200] = 3'b110;
        rom_memory[28201] = 3'b110;
        rom_memory[28202] = 3'b110;
        rom_memory[28203] = 3'b100;
        rom_memory[28204] = 3'b110;
        rom_memory[28205] = 3'b110;
        rom_memory[28206] = 3'b110;
        rom_memory[28207] = 3'b110;
        rom_memory[28208] = 3'b110;
        rom_memory[28209] = 3'b110;
        rom_memory[28210] = 3'b110;
        rom_memory[28211] = 3'b000;
        rom_memory[28212] = 3'b000;
        rom_memory[28213] = 3'b000;
        rom_memory[28214] = 3'b000;
        rom_memory[28215] = 3'b000;
        rom_memory[28216] = 3'b110;
        rom_memory[28217] = 3'b110;
        rom_memory[28218] = 3'b110;
        rom_memory[28219] = 3'b110;
        rom_memory[28220] = 3'b110;
        rom_memory[28221] = 3'b110;
        rom_memory[28222] = 3'b110;
        rom_memory[28223] = 3'b110;
        rom_memory[28224] = 3'b110;
        rom_memory[28225] = 3'b110;
        rom_memory[28226] = 3'b110;
        rom_memory[28227] = 3'b110;
        rom_memory[28228] = 3'b110;
        rom_memory[28229] = 3'b110;
        rom_memory[28230] = 3'b110;
        rom_memory[28231] = 3'b110;
        rom_memory[28232] = 3'b110;
        rom_memory[28233] = 3'b110;
        rom_memory[28234] = 3'b110;
        rom_memory[28235] = 3'b110;
        rom_memory[28236] = 3'b110;
        rom_memory[28237] = 3'b110;
        rom_memory[28238] = 3'b110;
        rom_memory[28239] = 3'b110;
        rom_memory[28240] = 3'b110;
        rom_memory[28241] = 3'b110;
        rom_memory[28242] = 3'b110;
        rom_memory[28243] = 3'b110;
        rom_memory[28244] = 3'b110;
        rom_memory[28245] = 3'b110;
        rom_memory[28246] = 3'b110;
        rom_memory[28247] = 3'b110;
        rom_memory[28248] = 3'b110;
        rom_memory[28249] = 3'b110;
        rom_memory[28250] = 3'b110;
        rom_memory[28251] = 3'b110;
        rom_memory[28252] = 3'b110;
        rom_memory[28253] = 3'b110;
        rom_memory[28254] = 3'b110;
        rom_memory[28255] = 3'b110;
        rom_memory[28256] = 3'b110;
        rom_memory[28257] = 3'b110;
        rom_memory[28258] = 3'b110;
        rom_memory[28259] = 3'b110;
        rom_memory[28260] = 3'b111;
        rom_memory[28261] = 3'b111;
        rom_memory[28262] = 3'b111;
        rom_memory[28263] = 3'b111;
        rom_memory[28264] = 3'b111;
        rom_memory[28265] = 3'b111;
        rom_memory[28266] = 3'b111;
        rom_memory[28267] = 3'b111;
        rom_memory[28268] = 3'b111;
        rom_memory[28269] = 3'b111;
        rom_memory[28270] = 3'b111;
        rom_memory[28271] = 3'b111;
        rom_memory[28272] = 3'b111;
        rom_memory[28273] = 3'b111;
        rom_memory[28274] = 3'b111;
        rom_memory[28275] = 3'b111;
        rom_memory[28276] = 3'b111;
        rom_memory[28277] = 3'b111;
        rom_memory[28278] = 3'b111;
        rom_memory[28279] = 3'b111;
        rom_memory[28280] = 3'b111;
        rom_memory[28281] = 3'b111;
        rom_memory[28282] = 3'b111;
        rom_memory[28283] = 3'b111;
        rom_memory[28284] = 3'b111;
        rom_memory[28285] = 3'b111;
        rom_memory[28286] = 3'b111;
        rom_memory[28287] = 3'b111;
        rom_memory[28288] = 3'b111;
        rom_memory[28289] = 3'b111;
        rom_memory[28290] = 3'b111;
        rom_memory[28291] = 3'b111;
        rom_memory[28292] = 3'b111;
        rom_memory[28293] = 3'b111;
        rom_memory[28294] = 3'b111;
        rom_memory[28295] = 3'b111;
        rom_memory[28296] = 3'b111;
        rom_memory[28297] = 3'b111;
        rom_memory[28298] = 3'b111;
        rom_memory[28299] = 3'b111;
        rom_memory[28300] = 3'b111;
        rom_memory[28301] = 3'b111;
        rom_memory[28302] = 3'b111;
        rom_memory[28303] = 3'b111;
        rom_memory[28304] = 3'b111;
        rom_memory[28305] = 3'b111;
        rom_memory[28306] = 3'b111;
        rom_memory[28307] = 3'b111;
        rom_memory[28308] = 3'b111;
        rom_memory[28309] = 3'b111;
        rom_memory[28310] = 3'b111;
        rom_memory[28311] = 3'b111;
        rom_memory[28312] = 3'b111;
        rom_memory[28313] = 3'b111;
        rom_memory[28314] = 3'b111;
        rom_memory[28315] = 3'b111;
        rom_memory[28316] = 3'b111;
        rom_memory[28317] = 3'b111;
        rom_memory[28318] = 3'b111;
        rom_memory[28319] = 3'b111;
        rom_memory[28320] = 3'b110;
        rom_memory[28321] = 3'b110;
        rom_memory[28322] = 3'b110;
        rom_memory[28323] = 3'b110;
        rom_memory[28324] = 3'b110;
        rom_memory[28325] = 3'b110;
        rom_memory[28326] = 3'b110;
        rom_memory[28327] = 3'b110;
        rom_memory[28328] = 3'b110;
        rom_memory[28329] = 3'b110;
        rom_memory[28330] = 3'b110;
        rom_memory[28331] = 3'b111;
        rom_memory[28332] = 3'b111;
        rom_memory[28333] = 3'b111;
        rom_memory[28334] = 3'b111;
        rom_memory[28335] = 3'b111;
        rom_memory[28336] = 3'b111;
        rom_memory[28337] = 3'b111;
        rom_memory[28338] = 3'b111;
        rom_memory[28339] = 3'b111;
        rom_memory[28340] = 3'b111;
        rom_memory[28341] = 3'b111;
        rom_memory[28342] = 3'b111;
        rom_memory[28343] = 3'b111;
        rom_memory[28344] = 3'b111;
        rom_memory[28345] = 3'b111;
        rom_memory[28346] = 3'b111;
        rom_memory[28347] = 3'b110;
        rom_memory[28348] = 3'b110;
        rom_memory[28349] = 3'b110;
        rom_memory[28350] = 3'b110;
        rom_memory[28351] = 3'b110;
        rom_memory[28352] = 3'b110;
        rom_memory[28353] = 3'b110;
        rom_memory[28354] = 3'b110;
        rom_memory[28355] = 3'b111;
        rom_memory[28356] = 3'b110;
        rom_memory[28357] = 3'b110;
        rom_memory[28358] = 3'b110;
        rom_memory[28359] = 3'b110;
        rom_memory[28360] = 3'b110;
        rom_memory[28361] = 3'b110;
        rom_memory[28362] = 3'b110;
        rom_memory[28363] = 3'b110;
        rom_memory[28364] = 3'b110;
        rom_memory[28365] = 3'b110;
        rom_memory[28366] = 3'b110;
        rom_memory[28367] = 3'b111;
        rom_memory[28368] = 3'b111;
        rom_memory[28369] = 3'b111;
        rom_memory[28370] = 3'b111;
        rom_memory[28371] = 3'b111;
        rom_memory[28372] = 3'b111;
        rom_memory[28373] = 3'b111;
        rom_memory[28374] = 3'b111;
        rom_memory[28375] = 3'b111;
        rom_memory[28376] = 3'b111;
        rom_memory[28377] = 3'b111;
        rom_memory[28378] = 3'b111;
        rom_memory[28379] = 3'b111;
        rom_memory[28380] = 3'b111;
        rom_memory[28381] = 3'b111;
        rom_memory[28382] = 3'b111;
        rom_memory[28383] = 3'b111;
        rom_memory[28384] = 3'b110;
        rom_memory[28385] = 3'b100;
        rom_memory[28386] = 3'b110;
        rom_memory[28387] = 3'b110;
        rom_memory[28388] = 3'b110;
        rom_memory[28389] = 3'b100;
        rom_memory[28390] = 3'b100;
        rom_memory[28391] = 3'b100;
        rom_memory[28392] = 3'b100;
        rom_memory[28393] = 3'b100;
        rom_memory[28394] = 3'b100;
        rom_memory[28395] = 3'b100;
        rom_memory[28396] = 3'b110;
        rom_memory[28397] = 3'b110;
        rom_memory[28398] = 3'b110;
        rom_memory[28399] = 3'b110;
        rom_memory[28400] = 3'b110;
        rom_memory[28401] = 3'b110;
        rom_memory[28402] = 3'b110;
        rom_memory[28403] = 3'b110;
        rom_memory[28404] = 3'b110;
        rom_memory[28405] = 3'b110;
        rom_memory[28406] = 3'b110;
        rom_memory[28407] = 3'b110;
        rom_memory[28408] = 3'b110;
        rom_memory[28409] = 3'b110;
        rom_memory[28410] = 3'b110;
        rom_memory[28411] = 3'b110;
        rom_memory[28412] = 3'b110;
        rom_memory[28413] = 3'b110;
        rom_memory[28414] = 3'b110;
        rom_memory[28415] = 3'b110;
        rom_memory[28416] = 3'b110;
        rom_memory[28417] = 3'b110;
        rom_memory[28418] = 3'b110;
        rom_memory[28419] = 3'b110;
        rom_memory[28420] = 3'b110;
        rom_memory[28421] = 3'b110;
        rom_memory[28422] = 3'b110;
        rom_memory[28423] = 3'b110;
        rom_memory[28424] = 3'b110;
        rom_memory[28425] = 3'b110;
        rom_memory[28426] = 3'b110;
        rom_memory[28427] = 3'b110;
        rom_memory[28428] = 3'b110;
        rom_memory[28429] = 3'b110;
        rom_memory[28430] = 3'b110;
        rom_memory[28431] = 3'b110;
        rom_memory[28432] = 3'b110;
        rom_memory[28433] = 3'b110;
        rom_memory[28434] = 3'b110;
        rom_memory[28435] = 3'b110;
        rom_memory[28436] = 3'b110;
        rom_memory[28437] = 3'b110;
        rom_memory[28438] = 3'b110;
        rom_memory[28439] = 3'b110;
        rom_memory[28440] = 3'b110;
        rom_memory[28441] = 3'b110;
        rom_memory[28442] = 3'b110;
        rom_memory[28443] = 3'b110;
        rom_memory[28444] = 3'b100;
        rom_memory[28445] = 3'b110;
        rom_memory[28446] = 3'b110;
        rom_memory[28447] = 3'b110;
        rom_memory[28448] = 3'b110;
        rom_memory[28449] = 3'b110;
        rom_memory[28450] = 3'b110;
        rom_memory[28451] = 3'b100;
        rom_memory[28452] = 3'b000;
        rom_memory[28453] = 3'b000;
        rom_memory[28454] = 3'b000;
        rom_memory[28455] = 3'b000;
        rom_memory[28456] = 3'b110;
        rom_memory[28457] = 3'b110;
        rom_memory[28458] = 3'b110;
        rom_memory[28459] = 3'b110;
        rom_memory[28460] = 3'b110;
        rom_memory[28461] = 3'b110;
        rom_memory[28462] = 3'b110;
        rom_memory[28463] = 3'b110;
        rom_memory[28464] = 3'b110;
        rom_memory[28465] = 3'b110;
        rom_memory[28466] = 3'b110;
        rom_memory[28467] = 3'b110;
        rom_memory[28468] = 3'b110;
        rom_memory[28469] = 3'b110;
        rom_memory[28470] = 3'b110;
        rom_memory[28471] = 3'b110;
        rom_memory[28472] = 3'b110;
        rom_memory[28473] = 3'b110;
        rom_memory[28474] = 3'b110;
        rom_memory[28475] = 3'b110;
        rom_memory[28476] = 3'b110;
        rom_memory[28477] = 3'b110;
        rom_memory[28478] = 3'b110;
        rom_memory[28479] = 3'b110;
        rom_memory[28480] = 3'b110;
        rom_memory[28481] = 3'b110;
        rom_memory[28482] = 3'b110;
        rom_memory[28483] = 3'b110;
        rom_memory[28484] = 3'b110;
        rom_memory[28485] = 3'b110;
        rom_memory[28486] = 3'b110;
        rom_memory[28487] = 3'b110;
        rom_memory[28488] = 3'b110;
        rom_memory[28489] = 3'b110;
        rom_memory[28490] = 3'b110;
        rom_memory[28491] = 3'b110;
        rom_memory[28492] = 3'b110;
        rom_memory[28493] = 3'b110;
        rom_memory[28494] = 3'b110;
        rom_memory[28495] = 3'b110;
        rom_memory[28496] = 3'b110;
        rom_memory[28497] = 3'b110;
        rom_memory[28498] = 3'b110;
        rom_memory[28499] = 3'b110;
        rom_memory[28500] = 3'b111;
        rom_memory[28501] = 3'b111;
        rom_memory[28502] = 3'b111;
        rom_memory[28503] = 3'b111;
        rom_memory[28504] = 3'b111;
        rom_memory[28505] = 3'b111;
        rom_memory[28506] = 3'b111;
        rom_memory[28507] = 3'b111;
        rom_memory[28508] = 3'b111;
        rom_memory[28509] = 3'b111;
        rom_memory[28510] = 3'b111;
        rom_memory[28511] = 3'b111;
        rom_memory[28512] = 3'b111;
        rom_memory[28513] = 3'b111;
        rom_memory[28514] = 3'b111;
        rom_memory[28515] = 3'b111;
        rom_memory[28516] = 3'b111;
        rom_memory[28517] = 3'b111;
        rom_memory[28518] = 3'b111;
        rom_memory[28519] = 3'b111;
        rom_memory[28520] = 3'b111;
        rom_memory[28521] = 3'b111;
        rom_memory[28522] = 3'b111;
        rom_memory[28523] = 3'b111;
        rom_memory[28524] = 3'b111;
        rom_memory[28525] = 3'b111;
        rom_memory[28526] = 3'b111;
        rom_memory[28527] = 3'b111;
        rom_memory[28528] = 3'b111;
        rom_memory[28529] = 3'b111;
        rom_memory[28530] = 3'b111;
        rom_memory[28531] = 3'b111;
        rom_memory[28532] = 3'b111;
        rom_memory[28533] = 3'b111;
        rom_memory[28534] = 3'b111;
        rom_memory[28535] = 3'b111;
        rom_memory[28536] = 3'b111;
        rom_memory[28537] = 3'b111;
        rom_memory[28538] = 3'b111;
        rom_memory[28539] = 3'b111;
        rom_memory[28540] = 3'b111;
        rom_memory[28541] = 3'b111;
        rom_memory[28542] = 3'b111;
        rom_memory[28543] = 3'b111;
        rom_memory[28544] = 3'b111;
        rom_memory[28545] = 3'b111;
        rom_memory[28546] = 3'b111;
        rom_memory[28547] = 3'b111;
        rom_memory[28548] = 3'b111;
        rom_memory[28549] = 3'b111;
        rom_memory[28550] = 3'b111;
        rom_memory[28551] = 3'b111;
        rom_memory[28552] = 3'b111;
        rom_memory[28553] = 3'b111;
        rom_memory[28554] = 3'b111;
        rom_memory[28555] = 3'b111;
        rom_memory[28556] = 3'b111;
        rom_memory[28557] = 3'b111;
        rom_memory[28558] = 3'b111;
        rom_memory[28559] = 3'b111;
        rom_memory[28560] = 3'b110;
        rom_memory[28561] = 3'b110;
        rom_memory[28562] = 3'b110;
        rom_memory[28563] = 3'b110;
        rom_memory[28564] = 3'b110;
        rom_memory[28565] = 3'b110;
        rom_memory[28566] = 3'b110;
        rom_memory[28567] = 3'b110;
        rom_memory[28568] = 3'b110;
        rom_memory[28569] = 3'b110;
        rom_memory[28570] = 3'b110;
        rom_memory[28571] = 3'b111;
        rom_memory[28572] = 3'b111;
        rom_memory[28573] = 3'b111;
        rom_memory[28574] = 3'b111;
        rom_memory[28575] = 3'b111;
        rom_memory[28576] = 3'b111;
        rom_memory[28577] = 3'b111;
        rom_memory[28578] = 3'b111;
        rom_memory[28579] = 3'b111;
        rom_memory[28580] = 3'b111;
        rom_memory[28581] = 3'b111;
        rom_memory[28582] = 3'b111;
        rom_memory[28583] = 3'b111;
        rom_memory[28584] = 3'b111;
        rom_memory[28585] = 3'b111;
        rom_memory[28586] = 3'b111;
        rom_memory[28587] = 3'b110;
        rom_memory[28588] = 3'b110;
        rom_memory[28589] = 3'b110;
        rom_memory[28590] = 3'b110;
        rom_memory[28591] = 3'b110;
        rom_memory[28592] = 3'b110;
        rom_memory[28593] = 3'b110;
        rom_memory[28594] = 3'b110;
        rom_memory[28595] = 3'b111;
        rom_memory[28596] = 3'b110;
        rom_memory[28597] = 3'b110;
        rom_memory[28598] = 3'b110;
        rom_memory[28599] = 3'b110;
        rom_memory[28600] = 3'b110;
        rom_memory[28601] = 3'b110;
        rom_memory[28602] = 3'b110;
        rom_memory[28603] = 3'b110;
        rom_memory[28604] = 3'b110;
        rom_memory[28605] = 3'b110;
        rom_memory[28606] = 3'b110;
        rom_memory[28607] = 3'b111;
        rom_memory[28608] = 3'b111;
        rom_memory[28609] = 3'b111;
        rom_memory[28610] = 3'b111;
        rom_memory[28611] = 3'b111;
        rom_memory[28612] = 3'b111;
        rom_memory[28613] = 3'b111;
        rom_memory[28614] = 3'b111;
        rom_memory[28615] = 3'b111;
        rom_memory[28616] = 3'b111;
        rom_memory[28617] = 3'b111;
        rom_memory[28618] = 3'b111;
        rom_memory[28619] = 3'b111;
        rom_memory[28620] = 3'b111;
        rom_memory[28621] = 3'b111;
        rom_memory[28622] = 3'b111;
        rom_memory[28623] = 3'b111;
        rom_memory[28624] = 3'b111;
        rom_memory[28625] = 3'b110;
        rom_memory[28626] = 3'b110;
        rom_memory[28627] = 3'b110;
        rom_memory[28628] = 3'b110;
        rom_memory[28629] = 3'b110;
        rom_memory[28630] = 3'b100;
        rom_memory[28631] = 3'b100;
        rom_memory[28632] = 3'b100;
        rom_memory[28633] = 3'b100;
        rom_memory[28634] = 3'b100;
        rom_memory[28635] = 3'b100;
        rom_memory[28636] = 3'b100;
        rom_memory[28637] = 3'b110;
        rom_memory[28638] = 3'b110;
        rom_memory[28639] = 3'b110;
        rom_memory[28640] = 3'b110;
        rom_memory[28641] = 3'b110;
        rom_memory[28642] = 3'b110;
        rom_memory[28643] = 3'b110;
        rom_memory[28644] = 3'b110;
        rom_memory[28645] = 3'b110;
        rom_memory[28646] = 3'b110;
        rom_memory[28647] = 3'b110;
        rom_memory[28648] = 3'b110;
        rom_memory[28649] = 3'b110;
        rom_memory[28650] = 3'b110;
        rom_memory[28651] = 3'b110;
        rom_memory[28652] = 3'b110;
        rom_memory[28653] = 3'b110;
        rom_memory[28654] = 3'b110;
        rom_memory[28655] = 3'b110;
        rom_memory[28656] = 3'b110;
        rom_memory[28657] = 3'b110;
        rom_memory[28658] = 3'b110;
        rom_memory[28659] = 3'b110;
        rom_memory[28660] = 3'b110;
        rom_memory[28661] = 3'b110;
        rom_memory[28662] = 3'b110;
        rom_memory[28663] = 3'b110;
        rom_memory[28664] = 3'b110;
        rom_memory[28665] = 3'b110;
        rom_memory[28666] = 3'b110;
        rom_memory[28667] = 3'b110;
        rom_memory[28668] = 3'b110;
        rom_memory[28669] = 3'b110;
        rom_memory[28670] = 3'b110;
        rom_memory[28671] = 3'b110;
        rom_memory[28672] = 3'b110;
        rom_memory[28673] = 3'b110;
        rom_memory[28674] = 3'b110;
        rom_memory[28675] = 3'b110;
        rom_memory[28676] = 3'b110;
        rom_memory[28677] = 3'b110;
        rom_memory[28678] = 3'b110;
        rom_memory[28679] = 3'b110;
        rom_memory[28680] = 3'b110;
        rom_memory[28681] = 3'b110;
        rom_memory[28682] = 3'b110;
        rom_memory[28683] = 3'b110;
        rom_memory[28684] = 3'b110;
        rom_memory[28685] = 3'b100;
        rom_memory[28686] = 3'b110;
        rom_memory[28687] = 3'b110;
        rom_memory[28688] = 3'b110;
        rom_memory[28689] = 3'b110;
        rom_memory[28690] = 3'b110;
        rom_memory[28691] = 3'b110;
        rom_memory[28692] = 3'b000;
        rom_memory[28693] = 3'b000;
        rom_memory[28694] = 3'b000;
        rom_memory[28695] = 3'b000;
        rom_memory[28696] = 3'b000;
        rom_memory[28697] = 3'b110;
        rom_memory[28698] = 3'b110;
        rom_memory[28699] = 3'b110;
        rom_memory[28700] = 3'b110;
        rom_memory[28701] = 3'b110;
        rom_memory[28702] = 3'b110;
        rom_memory[28703] = 3'b110;
        rom_memory[28704] = 3'b110;
        rom_memory[28705] = 3'b110;
        rom_memory[28706] = 3'b110;
        rom_memory[28707] = 3'b110;
        rom_memory[28708] = 3'b110;
        rom_memory[28709] = 3'b110;
        rom_memory[28710] = 3'b110;
        rom_memory[28711] = 3'b110;
        rom_memory[28712] = 3'b110;
        rom_memory[28713] = 3'b110;
        rom_memory[28714] = 3'b110;
        rom_memory[28715] = 3'b110;
        rom_memory[28716] = 3'b110;
        rom_memory[28717] = 3'b110;
        rom_memory[28718] = 3'b110;
        rom_memory[28719] = 3'b110;
        rom_memory[28720] = 3'b110;
        rom_memory[28721] = 3'b110;
        rom_memory[28722] = 3'b110;
        rom_memory[28723] = 3'b110;
        rom_memory[28724] = 3'b110;
        rom_memory[28725] = 3'b110;
        rom_memory[28726] = 3'b110;
        rom_memory[28727] = 3'b110;
        rom_memory[28728] = 3'b110;
        rom_memory[28729] = 3'b110;
        rom_memory[28730] = 3'b110;
        rom_memory[28731] = 3'b110;
        rom_memory[28732] = 3'b110;
        rom_memory[28733] = 3'b110;
        rom_memory[28734] = 3'b110;
        rom_memory[28735] = 3'b110;
        rom_memory[28736] = 3'b110;
        rom_memory[28737] = 3'b110;
        rom_memory[28738] = 3'b110;
        rom_memory[28739] = 3'b110;
        rom_memory[28740] = 3'b111;
        rom_memory[28741] = 3'b111;
        rom_memory[28742] = 3'b111;
        rom_memory[28743] = 3'b111;
        rom_memory[28744] = 3'b111;
        rom_memory[28745] = 3'b111;
        rom_memory[28746] = 3'b111;
        rom_memory[28747] = 3'b111;
        rom_memory[28748] = 3'b111;
        rom_memory[28749] = 3'b111;
        rom_memory[28750] = 3'b111;
        rom_memory[28751] = 3'b111;
        rom_memory[28752] = 3'b111;
        rom_memory[28753] = 3'b111;
        rom_memory[28754] = 3'b111;
        rom_memory[28755] = 3'b111;
        rom_memory[28756] = 3'b111;
        rom_memory[28757] = 3'b111;
        rom_memory[28758] = 3'b111;
        rom_memory[28759] = 3'b111;
        rom_memory[28760] = 3'b111;
        rom_memory[28761] = 3'b111;
        rom_memory[28762] = 3'b111;
        rom_memory[28763] = 3'b111;
        rom_memory[28764] = 3'b111;
        rom_memory[28765] = 3'b111;
        rom_memory[28766] = 3'b111;
        rom_memory[28767] = 3'b111;
        rom_memory[28768] = 3'b111;
        rom_memory[28769] = 3'b111;
        rom_memory[28770] = 3'b111;
        rom_memory[28771] = 3'b111;
        rom_memory[28772] = 3'b111;
        rom_memory[28773] = 3'b111;
        rom_memory[28774] = 3'b111;
        rom_memory[28775] = 3'b111;
        rom_memory[28776] = 3'b111;
        rom_memory[28777] = 3'b111;
        rom_memory[28778] = 3'b111;
        rom_memory[28779] = 3'b111;
        rom_memory[28780] = 3'b111;
        rom_memory[28781] = 3'b111;
        rom_memory[28782] = 3'b111;
        rom_memory[28783] = 3'b111;
        rom_memory[28784] = 3'b111;
        rom_memory[28785] = 3'b111;
        rom_memory[28786] = 3'b111;
        rom_memory[28787] = 3'b111;
        rom_memory[28788] = 3'b111;
        rom_memory[28789] = 3'b111;
        rom_memory[28790] = 3'b111;
        rom_memory[28791] = 3'b111;
        rom_memory[28792] = 3'b111;
        rom_memory[28793] = 3'b111;
        rom_memory[28794] = 3'b111;
        rom_memory[28795] = 3'b111;
        rom_memory[28796] = 3'b111;
        rom_memory[28797] = 3'b111;
        rom_memory[28798] = 3'b111;
        rom_memory[28799] = 3'b111;
        rom_memory[28800] = 3'b110;
        rom_memory[28801] = 3'b110;
        rom_memory[28802] = 3'b110;
        rom_memory[28803] = 3'b110;
        rom_memory[28804] = 3'b110;
        rom_memory[28805] = 3'b110;
        rom_memory[28806] = 3'b110;
        rom_memory[28807] = 3'b110;
        rom_memory[28808] = 3'b110;
        rom_memory[28809] = 3'b110;
        rom_memory[28810] = 3'b111;
        rom_memory[28811] = 3'b111;
        rom_memory[28812] = 3'b111;
        rom_memory[28813] = 3'b111;
        rom_memory[28814] = 3'b111;
        rom_memory[28815] = 3'b111;
        rom_memory[28816] = 3'b111;
        rom_memory[28817] = 3'b111;
        rom_memory[28818] = 3'b111;
        rom_memory[28819] = 3'b111;
        rom_memory[28820] = 3'b111;
        rom_memory[28821] = 3'b111;
        rom_memory[28822] = 3'b111;
        rom_memory[28823] = 3'b111;
        rom_memory[28824] = 3'b111;
        rom_memory[28825] = 3'b111;
        rom_memory[28826] = 3'b111;
        rom_memory[28827] = 3'b111;
        rom_memory[28828] = 3'b110;
        rom_memory[28829] = 3'b110;
        rom_memory[28830] = 3'b110;
        rom_memory[28831] = 3'b110;
        rom_memory[28832] = 3'b110;
        rom_memory[28833] = 3'b110;
        rom_memory[28834] = 3'b110;
        rom_memory[28835] = 3'b110;
        rom_memory[28836] = 3'b110;
        rom_memory[28837] = 3'b110;
        rom_memory[28838] = 3'b110;
        rom_memory[28839] = 3'b110;
        rom_memory[28840] = 3'b110;
        rom_memory[28841] = 3'b110;
        rom_memory[28842] = 3'b110;
        rom_memory[28843] = 3'b110;
        rom_memory[28844] = 3'b110;
        rom_memory[28845] = 3'b111;
        rom_memory[28846] = 3'b111;
        rom_memory[28847] = 3'b111;
        rom_memory[28848] = 3'b111;
        rom_memory[28849] = 3'b111;
        rom_memory[28850] = 3'b111;
        rom_memory[28851] = 3'b111;
        rom_memory[28852] = 3'b111;
        rom_memory[28853] = 3'b111;
        rom_memory[28854] = 3'b111;
        rom_memory[28855] = 3'b111;
        rom_memory[28856] = 3'b111;
        rom_memory[28857] = 3'b111;
        rom_memory[28858] = 3'b111;
        rom_memory[28859] = 3'b111;
        rom_memory[28860] = 3'b111;
        rom_memory[28861] = 3'b111;
        rom_memory[28862] = 3'b111;
        rom_memory[28863] = 3'b111;
        rom_memory[28864] = 3'b111;
        rom_memory[28865] = 3'b111;
        rom_memory[28866] = 3'b110;
        rom_memory[28867] = 3'b110;
        rom_memory[28868] = 3'b110;
        rom_memory[28869] = 3'b110;
        rom_memory[28870] = 3'b100;
        rom_memory[28871] = 3'b100;
        rom_memory[28872] = 3'b100;
        rom_memory[28873] = 3'b100;
        rom_memory[28874] = 3'b100;
        rom_memory[28875] = 3'b100;
        rom_memory[28876] = 3'b100;
        rom_memory[28877] = 3'b100;
        rom_memory[28878] = 3'b110;
        rom_memory[28879] = 3'b110;
        rom_memory[28880] = 3'b110;
        rom_memory[28881] = 3'b110;
        rom_memory[28882] = 3'b110;
        rom_memory[28883] = 3'b110;
        rom_memory[28884] = 3'b110;
        rom_memory[28885] = 3'b110;
        rom_memory[28886] = 3'b110;
        rom_memory[28887] = 3'b110;
        rom_memory[28888] = 3'b110;
        rom_memory[28889] = 3'b110;
        rom_memory[28890] = 3'b110;
        rom_memory[28891] = 3'b110;
        rom_memory[28892] = 3'b110;
        rom_memory[28893] = 3'b110;
        rom_memory[28894] = 3'b110;
        rom_memory[28895] = 3'b110;
        rom_memory[28896] = 3'b110;
        rom_memory[28897] = 3'b110;
        rom_memory[28898] = 3'b111;
        rom_memory[28899] = 3'b110;
        rom_memory[28900] = 3'b110;
        rom_memory[28901] = 3'b110;
        rom_memory[28902] = 3'b110;
        rom_memory[28903] = 3'b110;
        rom_memory[28904] = 3'b110;
        rom_memory[28905] = 3'b110;
        rom_memory[28906] = 3'b110;
        rom_memory[28907] = 3'b110;
        rom_memory[28908] = 3'b110;
        rom_memory[28909] = 3'b110;
        rom_memory[28910] = 3'b110;
        rom_memory[28911] = 3'b110;
        rom_memory[28912] = 3'b110;
        rom_memory[28913] = 3'b110;
        rom_memory[28914] = 3'b110;
        rom_memory[28915] = 3'b110;
        rom_memory[28916] = 3'b110;
        rom_memory[28917] = 3'b110;
        rom_memory[28918] = 3'b110;
        rom_memory[28919] = 3'b110;
        rom_memory[28920] = 3'b110;
        rom_memory[28921] = 3'b110;
        rom_memory[28922] = 3'b110;
        rom_memory[28923] = 3'b110;
        rom_memory[28924] = 3'b110;
        rom_memory[28925] = 3'b100;
        rom_memory[28926] = 3'b110;
        rom_memory[28927] = 3'b110;
        rom_memory[28928] = 3'b110;
        rom_memory[28929] = 3'b110;
        rom_memory[28930] = 3'b110;
        rom_memory[28931] = 3'b110;
        rom_memory[28932] = 3'b100;
        rom_memory[28933] = 3'b000;
        rom_memory[28934] = 3'b000;
        rom_memory[28935] = 3'b000;
        rom_memory[28936] = 3'b000;
        rom_memory[28937] = 3'b110;
        rom_memory[28938] = 3'b110;
        rom_memory[28939] = 3'b110;
        rom_memory[28940] = 3'b110;
        rom_memory[28941] = 3'b110;
        rom_memory[28942] = 3'b110;
        rom_memory[28943] = 3'b110;
        rom_memory[28944] = 3'b110;
        rom_memory[28945] = 3'b110;
        rom_memory[28946] = 3'b110;
        rom_memory[28947] = 3'b110;
        rom_memory[28948] = 3'b110;
        rom_memory[28949] = 3'b110;
        rom_memory[28950] = 3'b110;
        rom_memory[28951] = 3'b110;
        rom_memory[28952] = 3'b110;
        rom_memory[28953] = 3'b110;
        rom_memory[28954] = 3'b110;
        rom_memory[28955] = 3'b110;
        rom_memory[28956] = 3'b110;
        rom_memory[28957] = 3'b110;
        rom_memory[28958] = 3'b110;
        rom_memory[28959] = 3'b110;
        rom_memory[28960] = 3'b110;
        rom_memory[28961] = 3'b110;
        rom_memory[28962] = 3'b110;
        rom_memory[28963] = 3'b110;
        rom_memory[28964] = 3'b110;
        rom_memory[28965] = 3'b110;
        rom_memory[28966] = 3'b110;
        rom_memory[28967] = 3'b110;
        rom_memory[28968] = 3'b110;
        rom_memory[28969] = 3'b110;
        rom_memory[28970] = 3'b110;
        rom_memory[28971] = 3'b110;
        rom_memory[28972] = 3'b110;
        rom_memory[28973] = 3'b110;
        rom_memory[28974] = 3'b110;
        rom_memory[28975] = 3'b110;
        rom_memory[28976] = 3'b110;
        rom_memory[28977] = 3'b110;
        rom_memory[28978] = 3'b110;
        rom_memory[28979] = 3'b110;
        rom_memory[28980] = 3'b110;
        rom_memory[28981] = 3'b110;
        rom_memory[28982] = 3'b111;
        rom_memory[28983] = 3'b111;
        rom_memory[28984] = 3'b111;
        rom_memory[28985] = 3'b111;
        rom_memory[28986] = 3'b111;
        rom_memory[28987] = 3'b111;
        rom_memory[28988] = 3'b111;
        rom_memory[28989] = 3'b111;
        rom_memory[28990] = 3'b111;
        rom_memory[28991] = 3'b111;
        rom_memory[28992] = 3'b111;
        rom_memory[28993] = 3'b111;
        rom_memory[28994] = 3'b111;
        rom_memory[28995] = 3'b111;
        rom_memory[28996] = 3'b111;
        rom_memory[28997] = 3'b111;
        rom_memory[28998] = 3'b111;
        rom_memory[28999] = 3'b111;
        rom_memory[29000] = 3'b111;
        rom_memory[29001] = 3'b111;
        rom_memory[29002] = 3'b111;
        rom_memory[29003] = 3'b111;
        rom_memory[29004] = 3'b111;
        rom_memory[29005] = 3'b111;
        rom_memory[29006] = 3'b111;
        rom_memory[29007] = 3'b111;
        rom_memory[29008] = 3'b111;
        rom_memory[29009] = 3'b111;
        rom_memory[29010] = 3'b111;
        rom_memory[29011] = 3'b111;
        rom_memory[29012] = 3'b111;
        rom_memory[29013] = 3'b111;
        rom_memory[29014] = 3'b111;
        rom_memory[29015] = 3'b111;
        rom_memory[29016] = 3'b111;
        rom_memory[29017] = 3'b111;
        rom_memory[29018] = 3'b111;
        rom_memory[29019] = 3'b111;
        rom_memory[29020] = 3'b111;
        rom_memory[29021] = 3'b111;
        rom_memory[29022] = 3'b111;
        rom_memory[29023] = 3'b111;
        rom_memory[29024] = 3'b111;
        rom_memory[29025] = 3'b111;
        rom_memory[29026] = 3'b111;
        rom_memory[29027] = 3'b111;
        rom_memory[29028] = 3'b111;
        rom_memory[29029] = 3'b111;
        rom_memory[29030] = 3'b111;
        rom_memory[29031] = 3'b111;
        rom_memory[29032] = 3'b111;
        rom_memory[29033] = 3'b111;
        rom_memory[29034] = 3'b111;
        rom_memory[29035] = 3'b111;
        rom_memory[29036] = 3'b111;
        rom_memory[29037] = 3'b111;
        rom_memory[29038] = 3'b111;
        rom_memory[29039] = 3'b111;
        rom_memory[29040] = 3'b110;
        rom_memory[29041] = 3'b110;
        rom_memory[29042] = 3'b110;
        rom_memory[29043] = 3'b110;
        rom_memory[29044] = 3'b110;
        rom_memory[29045] = 3'b110;
        rom_memory[29046] = 3'b110;
        rom_memory[29047] = 3'b110;
        rom_memory[29048] = 3'b110;
        rom_memory[29049] = 3'b110;
        rom_memory[29050] = 3'b111;
        rom_memory[29051] = 3'b111;
        rom_memory[29052] = 3'b111;
        rom_memory[29053] = 3'b111;
        rom_memory[29054] = 3'b111;
        rom_memory[29055] = 3'b111;
        rom_memory[29056] = 3'b111;
        rom_memory[29057] = 3'b111;
        rom_memory[29058] = 3'b111;
        rom_memory[29059] = 3'b111;
        rom_memory[29060] = 3'b111;
        rom_memory[29061] = 3'b111;
        rom_memory[29062] = 3'b111;
        rom_memory[29063] = 3'b111;
        rom_memory[29064] = 3'b111;
        rom_memory[29065] = 3'b111;
        rom_memory[29066] = 3'b111;
        rom_memory[29067] = 3'b111;
        rom_memory[29068] = 3'b110;
        rom_memory[29069] = 3'b110;
        rom_memory[29070] = 3'b110;
        rom_memory[29071] = 3'b110;
        rom_memory[29072] = 3'b111;
        rom_memory[29073] = 3'b110;
        rom_memory[29074] = 3'b110;
        rom_memory[29075] = 3'b110;
        rom_memory[29076] = 3'b110;
        rom_memory[29077] = 3'b110;
        rom_memory[29078] = 3'b110;
        rom_memory[29079] = 3'b110;
        rom_memory[29080] = 3'b110;
        rom_memory[29081] = 3'b110;
        rom_memory[29082] = 3'b110;
        rom_memory[29083] = 3'b110;
        rom_memory[29084] = 3'b110;
        rom_memory[29085] = 3'b111;
        rom_memory[29086] = 3'b111;
        rom_memory[29087] = 3'b111;
        rom_memory[29088] = 3'b111;
        rom_memory[29089] = 3'b111;
        rom_memory[29090] = 3'b111;
        rom_memory[29091] = 3'b111;
        rom_memory[29092] = 3'b111;
        rom_memory[29093] = 3'b111;
        rom_memory[29094] = 3'b111;
        rom_memory[29095] = 3'b111;
        rom_memory[29096] = 3'b111;
        rom_memory[29097] = 3'b111;
        rom_memory[29098] = 3'b111;
        rom_memory[29099] = 3'b111;
        rom_memory[29100] = 3'b111;
        rom_memory[29101] = 3'b111;
        rom_memory[29102] = 3'b111;
        rom_memory[29103] = 3'b111;
        rom_memory[29104] = 3'b111;
        rom_memory[29105] = 3'b111;
        rom_memory[29106] = 3'b111;
        rom_memory[29107] = 3'b110;
        rom_memory[29108] = 3'b110;
        rom_memory[29109] = 3'b110;
        rom_memory[29110] = 3'b110;
        rom_memory[29111] = 3'b100;
        rom_memory[29112] = 3'b100;
        rom_memory[29113] = 3'b100;
        rom_memory[29114] = 3'b100;
        rom_memory[29115] = 3'b100;
        rom_memory[29116] = 3'b100;
        rom_memory[29117] = 3'b100;
        rom_memory[29118] = 3'b110;
        rom_memory[29119] = 3'b110;
        rom_memory[29120] = 3'b110;
        rom_memory[29121] = 3'b110;
        rom_memory[29122] = 3'b110;
        rom_memory[29123] = 3'b110;
        rom_memory[29124] = 3'b110;
        rom_memory[29125] = 3'b110;
        rom_memory[29126] = 3'b110;
        rom_memory[29127] = 3'b110;
        rom_memory[29128] = 3'b110;
        rom_memory[29129] = 3'b110;
        rom_memory[29130] = 3'b110;
        rom_memory[29131] = 3'b110;
        rom_memory[29132] = 3'b110;
        rom_memory[29133] = 3'b110;
        rom_memory[29134] = 3'b110;
        rom_memory[29135] = 3'b110;
        rom_memory[29136] = 3'b110;
        rom_memory[29137] = 3'b111;
        rom_memory[29138] = 3'b111;
        rom_memory[29139] = 3'b110;
        rom_memory[29140] = 3'b110;
        rom_memory[29141] = 3'b110;
        rom_memory[29142] = 3'b110;
        rom_memory[29143] = 3'b110;
        rom_memory[29144] = 3'b110;
        rom_memory[29145] = 3'b110;
        rom_memory[29146] = 3'b110;
        rom_memory[29147] = 3'b110;
        rom_memory[29148] = 3'b110;
        rom_memory[29149] = 3'b110;
        rom_memory[29150] = 3'b110;
        rom_memory[29151] = 3'b110;
        rom_memory[29152] = 3'b110;
        rom_memory[29153] = 3'b110;
        rom_memory[29154] = 3'b110;
        rom_memory[29155] = 3'b110;
        rom_memory[29156] = 3'b110;
        rom_memory[29157] = 3'b110;
        rom_memory[29158] = 3'b110;
        rom_memory[29159] = 3'b110;
        rom_memory[29160] = 3'b110;
        rom_memory[29161] = 3'b110;
        rom_memory[29162] = 3'b110;
        rom_memory[29163] = 3'b110;
        rom_memory[29164] = 3'b110;
        rom_memory[29165] = 3'b110;
        rom_memory[29166] = 3'b100;
        rom_memory[29167] = 3'b110;
        rom_memory[29168] = 3'b110;
        rom_memory[29169] = 3'b110;
        rom_memory[29170] = 3'b110;
        rom_memory[29171] = 3'b110;
        rom_memory[29172] = 3'b110;
        rom_memory[29173] = 3'b100;
        rom_memory[29174] = 3'b000;
        rom_memory[29175] = 3'b111;
        rom_memory[29176] = 3'b111;
        rom_memory[29177] = 3'b110;
        rom_memory[29178] = 3'b110;
        rom_memory[29179] = 3'b110;
        rom_memory[29180] = 3'b110;
        rom_memory[29181] = 3'b110;
        rom_memory[29182] = 3'b110;
        rom_memory[29183] = 3'b110;
        rom_memory[29184] = 3'b110;
        rom_memory[29185] = 3'b110;
        rom_memory[29186] = 3'b110;
        rom_memory[29187] = 3'b110;
        rom_memory[29188] = 3'b110;
        rom_memory[29189] = 3'b110;
        rom_memory[29190] = 3'b110;
        rom_memory[29191] = 3'b110;
        rom_memory[29192] = 3'b110;
        rom_memory[29193] = 3'b110;
        rom_memory[29194] = 3'b110;
        rom_memory[29195] = 3'b110;
        rom_memory[29196] = 3'b110;
        rom_memory[29197] = 3'b110;
        rom_memory[29198] = 3'b110;
        rom_memory[29199] = 3'b110;
        rom_memory[29200] = 3'b110;
        rom_memory[29201] = 3'b110;
        rom_memory[29202] = 3'b110;
        rom_memory[29203] = 3'b110;
        rom_memory[29204] = 3'b110;
        rom_memory[29205] = 3'b110;
        rom_memory[29206] = 3'b110;
        rom_memory[29207] = 3'b110;
        rom_memory[29208] = 3'b110;
        rom_memory[29209] = 3'b110;
        rom_memory[29210] = 3'b110;
        rom_memory[29211] = 3'b110;
        rom_memory[29212] = 3'b110;
        rom_memory[29213] = 3'b110;
        rom_memory[29214] = 3'b110;
        rom_memory[29215] = 3'b110;
        rom_memory[29216] = 3'b110;
        rom_memory[29217] = 3'b110;
        rom_memory[29218] = 3'b110;
        rom_memory[29219] = 3'b110;
        rom_memory[29220] = 3'b110;
        rom_memory[29221] = 3'b110;
        rom_memory[29222] = 3'b111;
        rom_memory[29223] = 3'b111;
        rom_memory[29224] = 3'b111;
        rom_memory[29225] = 3'b111;
        rom_memory[29226] = 3'b111;
        rom_memory[29227] = 3'b111;
        rom_memory[29228] = 3'b111;
        rom_memory[29229] = 3'b111;
        rom_memory[29230] = 3'b111;
        rom_memory[29231] = 3'b111;
        rom_memory[29232] = 3'b111;
        rom_memory[29233] = 3'b111;
        rom_memory[29234] = 3'b111;
        rom_memory[29235] = 3'b111;
        rom_memory[29236] = 3'b111;
        rom_memory[29237] = 3'b111;
        rom_memory[29238] = 3'b111;
        rom_memory[29239] = 3'b111;
        rom_memory[29240] = 3'b111;
        rom_memory[29241] = 3'b111;
        rom_memory[29242] = 3'b111;
        rom_memory[29243] = 3'b111;
        rom_memory[29244] = 3'b111;
        rom_memory[29245] = 3'b111;
        rom_memory[29246] = 3'b111;
        rom_memory[29247] = 3'b111;
        rom_memory[29248] = 3'b111;
        rom_memory[29249] = 3'b111;
        rom_memory[29250] = 3'b111;
        rom_memory[29251] = 3'b111;
        rom_memory[29252] = 3'b111;
        rom_memory[29253] = 3'b111;
        rom_memory[29254] = 3'b111;
        rom_memory[29255] = 3'b111;
        rom_memory[29256] = 3'b111;
        rom_memory[29257] = 3'b111;
        rom_memory[29258] = 3'b111;
        rom_memory[29259] = 3'b111;
        rom_memory[29260] = 3'b111;
        rom_memory[29261] = 3'b111;
        rom_memory[29262] = 3'b111;
        rom_memory[29263] = 3'b111;
        rom_memory[29264] = 3'b111;
        rom_memory[29265] = 3'b111;
        rom_memory[29266] = 3'b111;
        rom_memory[29267] = 3'b111;
        rom_memory[29268] = 3'b111;
        rom_memory[29269] = 3'b111;
        rom_memory[29270] = 3'b111;
        rom_memory[29271] = 3'b111;
        rom_memory[29272] = 3'b111;
        rom_memory[29273] = 3'b111;
        rom_memory[29274] = 3'b111;
        rom_memory[29275] = 3'b111;
        rom_memory[29276] = 3'b111;
        rom_memory[29277] = 3'b111;
        rom_memory[29278] = 3'b111;
        rom_memory[29279] = 3'b111;
        rom_memory[29280] = 3'b110;
        rom_memory[29281] = 3'b110;
        rom_memory[29282] = 3'b110;
        rom_memory[29283] = 3'b110;
        rom_memory[29284] = 3'b110;
        rom_memory[29285] = 3'b110;
        rom_memory[29286] = 3'b110;
        rom_memory[29287] = 3'b110;
        rom_memory[29288] = 3'b110;
        rom_memory[29289] = 3'b110;
        rom_memory[29290] = 3'b111;
        rom_memory[29291] = 3'b111;
        rom_memory[29292] = 3'b111;
        rom_memory[29293] = 3'b111;
        rom_memory[29294] = 3'b111;
        rom_memory[29295] = 3'b111;
        rom_memory[29296] = 3'b111;
        rom_memory[29297] = 3'b111;
        rom_memory[29298] = 3'b111;
        rom_memory[29299] = 3'b111;
        rom_memory[29300] = 3'b111;
        rom_memory[29301] = 3'b111;
        rom_memory[29302] = 3'b111;
        rom_memory[29303] = 3'b111;
        rom_memory[29304] = 3'b111;
        rom_memory[29305] = 3'b111;
        rom_memory[29306] = 3'b111;
        rom_memory[29307] = 3'b111;
        rom_memory[29308] = 3'b111;
        rom_memory[29309] = 3'b110;
        rom_memory[29310] = 3'b110;
        rom_memory[29311] = 3'b110;
        rom_memory[29312] = 3'b110;
        rom_memory[29313] = 3'b110;
        rom_memory[29314] = 3'b110;
        rom_memory[29315] = 3'b110;
        rom_memory[29316] = 3'b110;
        rom_memory[29317] = 3'b110;
        rom_memory[29318] = 3'b110;
        rom_memory[29319] = 3'b110;
        rom_memory[29320] = 3'b110;
        rom_memory[29321] = 3'b110;
        rom_memory[29322] = 3'b110;
        rom_memory[29323] = 3'b110;
        rom_memory[29324] = 3'b110;
        rom_memory[29325] = 3'b111;
        rom_memory[29326] = 3'b111;
        rom_memory[29327] = 3'b111;
        rom_memory[29328] = 3'b111;
        rom_memory[29329] = 3'b111;
        rom_memory[29330] = 3'b111;
        rom_memory[29331] = 3'b111;
        rom_memory[29332] = 3'b111;
        rom_memory[29333] = 3'b111;
        rom_memory[29334] = 3'b111;
        rom_memory[29335] = 3'b111;
        rom_memory[29336] = 3'b111;
        rom_memory[29337] = 3'b111;
        rom_memory[29338] = 3'b111;
        rom_memory[29339] = 3'b111;
        rom_memory[29340] = 3'b111;
        rom_memory[29341] = 3'b111;
        rom_memory[29342] = 3'b111;
        rom_memory[29343] = 3'b111;
        rom_memory[29344] = 3'b111;
        rom_memory[29345] = 3'b111;
        rom_memory[29346] = 3'b111;
        rom_memory[29347] = 3'b111;
        rom_memory[29348] = 3'b111;
        rom_memory[29349] = 3'b110;
        rom_memory[29350] = 3'b110;
        rom_memory[29351] = 3'b110;
        rom_memory[29352] = 3'b100;
        rom_memory[29353] = 3'b100;
        rom_memory[29354] = 3'b100;
        rom_memory[29355] = 3'b100;
        rom_memory[29356] = 3'b100;
        rom_memory[29357] = 3'b100;
        rom_memory[29358] = 3'b100;
        rom_memory[29359] = 3'b100;
        rom_memory[29360] = 3'b100;
        rom_memory[29361] = 3'b100;
        rom_memory[29362] = 3'b100;
        rom_memory[29363] = 3'b110;
        rom_memory[29364] = 3'b110;
        rom_memory[29365] = 3'b110;
        rom_memory[29366] = 3'b110;
        rom_memory[29367] = 3'b110;
        rom_memory[29368] = 3'b110;
        rom_memory[29369] = 3'b110;
        rom_memory[29370] = 3'b110;
        rom_memory[29371] = 3'b110;
        rom_memory[29372] = 3'b110;
        rom_memory[29373] = 3'b111;
        rom_memory[29374] = 3'b110;
        rom_memory[29375] = 3'b110;
        rom_memory[29376] = 3'b111;
        rom_memory[29377] = 3'b111;
        rom_memory[29378] = 3'b110;
        rom_memory[29379] = 3'b110;
        rom_memory[29380] = 3'b110;
        rom_memory[29381] = 3'b110;
        rom_memory[29382] = 3'b110;
        rom_memory[29383] = 3'b110;
        rom_memory[29384] = 3'b110;
        rom_memory[29385] = 3'b110;
        rom_memory[29386] = 3'b110;
        rom_memory[29387] = 3'b110;
        rom_memory[29388] = 3'b110;
        rom_memory[29389] = 3'b110;
        rom_memory[29390] = 3'b110;
        rom_memory[29391] = 3'b110;
        rom_memory[29392] = 3'b110;
        rom_memory[29393] = 3'b110;
        rom_memory[29394] = 3'b110;
        rom_memory[29395] = 3'b100;
        rom_memory[29396] = 3'b100;
        rom_memory[29397] = 3'b110;
        rom_memory[29398] = 3'b100;
        rom_memory[29399] = 3'b100;
        rom_memory[29400] = 3'b110;
        rom_memory[29401] = 3'b110;
        rom_memory[29402] = 3'b110;
        rom_memory[29403] = 3'b110;
        rom_memory[29404] = 3'b110;
        rom_memory[29405] = 3'b110;
        rom_memory[29406] = 3'b100;
        rom_memory[29407] = 3'b100;
        rom_memory[29408] = 3'b110;
        rom_memory[29409] = 3'b110;
        rom_memory[29410] = 3'b110;
        rom_memory[29411] = 3'b110;
        rom_memory[29412] = 3'b110;
        rom_memory[29413] = 3'b110;
        rom_memory[29414] = 3'b100;
        rom_memory[29415] = 3'b111;
        rom_memory[29416] = 3'b111;
        rom_memory[29417] = 3'b110;
        rom_memory[29418] = 3'b110;
        rom_memory[29419] = 3'b110;
        rom_memory[29420] = 3'b110;
        rom_memory[29421] = 3'b110;
        rom_memory[29422] = 3'b110;
        rom_memory[29423] = 3'b110;
        rom_memory[29424] = 3'b110;
        rom_memory[29425] = 3'b110;
        rom_memory[29426] = 3'b110;
        rom_memory[29427] = 3'b110;
        rom_memory[29428] = 3'b110;
        rom_memory[29429] = 3'b110;
        rom_memory[29430] = 3'b110;
        rom_memory[29431] = 3'b110;
        rom_memory[29432] = 3'b110;
        rom_memory[29433] = 3'b110;
        rom_memory[29434] = 3'b110;
        rom_memory[29435] = 3'b110;
        rom_memory[29436] = 3'b110;
        rom_memory[29437] = 3'b110;
        rom_memory[29438] = 3'b110;
        rom_memory[29439] = 3'b110;
        rom_memory[29440] = 3'b110;
        rom_memory[29441] = 3'b110;
        rom_memory[29442] = 3'b110;
        rom_memory[29443] = 3'b110;
        rom_memory[29444] = 3'b110;
        rom_memory[29445] = 3'b110;
        rom_memory[29446] = 3'b110;
        rom_memory[29447] = 3'b110;
        rom_memory[29448] = 3'b110;
        rom_memory[29449] = 3'b110;
        rom_memory[29450] = 3'b110;
        rom_memory[29451] = 3'b110;
        rom_memory[29452] = 3'b110;
        rom_memory[29453] = 3'b110;
        rom_memory[29454] = 3'b110;
        rom_memory[29455] = 3'b110;
        rom_memory[29456] = 3'b110;
        rom_memory[29457] = 3'b110;
        rom_memory[29458] = 3'b110;
        rom_memory[29459] = 3'b110;
        rom_memory[29460] = 3'b110;
        rom_memory[29461] = 3'b110;
        rom_memory[29462] = 3'b111;
        rom_memory[29463] = 3'b111;
        rom_memory[29464] = 3'b111;
        rom_memory[29465] = 3'b111;
        rom_memory[29466] = 3'b111;
        rom_memory[29467] = 3'b111;
        rom_memory[29468] = 3'b111;
        rom_memory[29469] = 3'b111;
        rom_memory[29470] = 3'b111;
        rom_memory[29471] = 3'b111;
        rom_memory[29472] = 3'b111;
        rom_memory[29473] = 3'b111;
        rom_memory[29474] = 3'b111;
        rom_memory[29475] = 3'b111;
        rom_memory[29476] = 3'b111;
        rom_memory[29477] = 3'b111;
        rom_memory[29478] = 3'b111;
        rom_memory[29479] = 3'b111;
        rom_memory[29480] = 3'b111;
        rom_memory[29481] = 3'b111;
        rom_memory[29482] = 3'b111;
        rom_memory[29483] = 3'b111;
        rom_memory[29484] = 3'b111;
        rom_memory[29485] = 3'b111;
        rom_memory[29486] = 3'b111;
        rom_memory[29487] = 3'b111;
        rom_memory[29488] = 3'b111;
        rom_memory[29489] = 3'b111;
        rom_memory[29490] = 3'b111;
        rom_memory[29491] = 3'b111;
        rom_memory[29492] = 3'b111;
        rom_memory[29493] = 3'b111;
        rom_memory[29494] = 3'b111;
        rom_memory[29495] = 3'b111;
        rom_memory[29496] = 3'b111;
        rom_memory[29497] = 3'b111;
        rom_memory[29498] = 3'b111;
        rom_memory[29499] = 3'b111;
        rom_memory[29500] = 3'b111;
        rom_memory[29501] = 3'b111;
        rom_memory[29502] = 3'b111;
        rom_memory[29503] = 3'b111;
        rom_memory[29504] = 3'b111;
        rom_memory[29505] = 3'b111;
        rom_memory[29506] = 3'b111;
        rom_memory[29507] = 3'b111;
        rom_memory[29508] = 3'b111;
        rom_memory[29509] = 3'b111;
        rom_memory[29510] = 3'b111;
        rom_memory[29511] = 3'b111;
        rom_memory[29512] = 3'b111;
        rom_memory[29513] = 3'b111;
        rom_memory[29514] = 3'b111;
        rom_memory[29515] = 3'b111;
        rom_memory[29516] = 3'b111;
        rom_memory[29517] = 3'b111;
        rom_memory[29518] = 3'b111;
        rom_memory[29519] = 3'b111;
        rom_memory[29520] = 3'b110;
        rom_memory[29521] = 3'b110;
        rom_memory[29522] = 3'b110;
        rom_memory[29523] = 3'b110;
        rom_memory[29524] = 3'b110;
        rom_memory[29525] = 3'b110;
        rom_memory[29526] = 3'b110;
        rom_memory[29527] = 3'b110;
        rom_memory[29528] = 3'b110;
        rom_memory[29529] = 3'b110;
        rom_memory[29530] = 3'b110;
        rom_memory[29531] = 3'b111;
        rom_memory[29532] = 3'b111;
        rom_memory[29533] = 3'b111;
        rom_memory[29534] = 3'b111;
        rom_memory[29535] = 3'b111;
        rom_memory[29536] = 3'b111;
        rom_memory[29537] = 3'b111;
        rom_memory[29538] = 3'b111;
        rom_memory[29539] = 3'b111;
        rom_memory[29540] = 3'b111;
        rom_memory[29541] = 3'b111;
        rom_memory[29542] = 3'b111;
        rom_memory[29543] = 3'b111;
        rom_memory[29544] = 3'b111;
        rom_memory[29545] = 3'b111;
        rom_memory[29546] = 3'b111;
        rom_memory[29547] = 3'b111;
        rom_memory[29548] = 3'b111;
        rom_memory[29549] = 3'b110;
        rom_memory[29550] = 3'b110;
        rom_memory[29551] = 3'b110;
        rom_memory[29552] = 3'b110;
        rom_memory[29553] = 3'b110;
        rom_memory[29554] = 3'b110;
        rom_memory[29555] = 3'b110;
        rom_memory[29556] = 3'b110;
        rom_memory[29557] = 3'b110;
        rom_memory[29558] = 3'b110;
        rom_memory[29559] = 3'b110;
        rom_memory[29560] = 3'b110;
        rom_memory[29561] = 3'b110;
        rom_memory[29562] = 3'b110;
        rom_memory[29563] = 3'b110;
        rom_memory[29564] = 3'b110;
        rom_memory[29565] = 3'b111;
        rom_memory[29566] = 3'b111;
        rom_memory[29567] = 3'b111;
        rom_memory[29568] = 3'b111;
        rom_memory[29569] = 3'b111;
        rom_memory[29570] = 3'b111;
        rom_memory[29571] = 3'b111;
        rom_memory[29572] = 3'b111;
        rom_memory[29573] = 3'b111;
        rom_memory[29574] = 3'b111;
        rom_memory[29575] = 3'b111;
        rom_memory[29576] = 3'b111;
        rom_memory[29577] = 3'b111;
        rom_memory[29578] = 3'b111;
        rom_memory[29579] = 3'b111;
        rom_memory[29580] = 3'b111;
        rom_memory[29581] = 3'b111;
        rom_memory[29582] = 3'b111;
        rom_memory[29583] = 3'b111;
        rom_memory[29584] = 3'b111;
        rom_memory[29585] = 3'b111;
        rom_memory[29586] = 3'b111;
        rom_memory[29587] = 3'b111;
        rom_memory[29588] = 3'b111;
        rom_memory[29589] = 3'b111;
        rom_memory[29590] = 3'b110;
        rom_memory[29591] = 3'b110;
        rom_memory[29592] = 3'b110;
        rom_memory[29593] = 3'b100;
        rom_memory[29594] = 3'b100;
        rom_memory[29595] = 3'b100;
        rom_memory[29596] = 3'b100;
        rom_memory[29597] = 3'b100;
        rom_memory[29598] = 3'b100;
        rom_memory[29599] = 3'b100;
        rom_memory[29600] = 3'b100;
        rom_memory[29601] = 3'b100;
        rom_memory[29602] = 3'b100;
        rom_memory[29603] = 3'b100;
        rom_memory[29604] = 3'b100;
        rom_memory[29605] = 3'b110;
        rom_memory[29606] = 3'b110;
        rom_memory[29607] = 3'b110;
        rom_memory[29608] = 3'b110;
        rom_memory[29609] = 3'b110;
        rom_memory[29610] = 3'b110;
        rom_memory[29611] = 3'b110;
        rom_memory[29612] = 3'b110;
        rom_memory[29613] = 3'b111;
        rom_memory[29614] = 3'b110;
        rom_memory[29615] = 3'b111;
        rom_memory[29616] = 3'b111;
        rom_memory[29617] = 3'b111;
        rom_memory[29618] = 3'b110;
        rom_memory[29619] = 3'b110;
        rom_memory[29620] = 3'b110;
        rom_memory[29621] = 3'b110;
        rom_memory[29622] = 3'b110;
        rom_memory[29623] = 3'b110;
        rom_memory[29624] = 3'b110;
        rom_memory[29625] = 3'b110;
        rom_memory[29626] = 3'b110;
        rom_memory[29627] = 3'b110;
        rom_memory[29628] = 3'b110;
        rom_memory[29629] = 3'b110;
        rom_memory[29630] = 3'b110;
        rom_memory[29631] = 3'b110;
        rom_memory[29632] = 3'b110;
        rom_memory[29633] = 3'b110;
        rom_memory[29634] = 3'b100;
        rom_memory[29635] = 3'b100;
        rom_memory[29636] = 3'b100;
        rom_memory[29637] = 3'b100;
        rom_memory[29638] = 3'b100;
        rom_memory[29639] = 3'b110;
        rom_memory[29640] = 3'b110;
        rom_memory[29641] = 3'b110;
        rom_memory[29642] = 3'b110;
        rom_memory[29643] = 3'b110;
        rom_memory[29644] = 3'b110;
        rom_memory[29645] = 3'b110;
        rom_memory[29646] = 3'b110;
        rom_memory[29647] = 3'b100;
        rom_memory[29648] = 3'b100;
        rom_memory[29649] = 3'b110;
        rom_memory[29650] = 3'b110;
        rom_memory[29651] = 3'b110;
        rom_memory[29652] = 3'b110;
        rom_memory[29653] = 3'b110;
        rom_memory[29654] = 3'b110;
        rom_memory[29655] = 3'b100;
        rom_memory[29656] = 3'b111;
        rom_memory[29657] = 3'b111;
        rom_memory[29658] = 3'b110;
        rom_memory[29659] = 3'b110;
        rom_memory[29660] = 3'b110;
        rom_memory[29661] = 3'b110;
        rom_memory[29662] = 3'b110;
        rom_memory[29663] = 3'b110;
        rom_memory[29664] = 3'b110;
        rom_memory[29665] = 3'b110;
        rom_memory[29666] = 3'b110;
        rom_memory[29667] = 3'b110;
        rom_memory[29668] = 3'b110;
        rom_memory[29669] = 3'b110;
        rom_memory[29670] = 3'b110;
        rom_memory[29671] = 3'b110;
        rom_memory[29672] = 3'b110;
        rom_memory[29673] = 3'b110;
        rom_memory[29674] = 3'b110;
        rom_memory[29675] = 3'b110;
        rom_memory[29676] = 3'b110;
        rom_memory[29677] = 3'b110;
        rom_memory[29678] = 3'b110;
        rom_memory[29679] = 3'b110;
        rom_memory[29680] = 3'b110;
        rom_memory[29681] = 3'b110;
        rom_memory[29682] = 3'b110;
        rom_memory[29683] = 3'b110;
        rom_memory[29684] = 3'b110;
        rom_memory[29685] = 3'b110;
        rom_memory[29686] = 3'b110;
        rom_memory[29687] = 3'b110;
        rom_memory[29688] = 3'b110;
        rom_memory[29689] = 3'b110;
        rom_memory[29690] = 3'b110;
        rom_memory[29691] = 3'b110;
        rom_memory[29692] = 3'b110;
        rom_memory[29693] = 3'b110;
        rom_memory[29694] = 3'b110;
        rom_memory[29695] = 3'b110;
        rom_memory[29696] = 3'b110;
        rom_memory[29697] = 3'b110;
        rom_memory[29698] = 3'b110;
        rom_memory[29699] = 3'b110;
        rom_memory[29700] = 3'b110;
        rom_memory[29701] = 3'b110;
        rom_memory[29702] = 3'b111;
        rom_memory[29703] = 3'b111;
        rom_memory[29704] = 3'b111;
        rom_memory[29705] = 3'b111;
        rom_memory[29706] = 3'b111;
        rom_memory[29707] = 3'b111;
        rom_memory[29708] = 3'b111;
        rom_memory[29709] = 3'b111;
        rom_memory[29710] = 3'b111;
        rom_memory[29711] = 3'b111;
        rom_memory[29712] = 3'b111;
        rom_memory[29713] = 3'b111;
        rom_memory[29714] = 3'b111;
        rom_memory[29715] = 3'b111;
        rom_memory[29716] = 3'b111;
        rom_memory[29717] = 3'b111;
        rom_memory[29718] = 3'b111;
        rom_memory[29719] = 3'b111;
        rom_memory[29720] = 3'b111;
        rom_memory[29721] = 3'b111;
        rom_memory[29722] = 3'b111;
        rom_memory[29723] = 3'b111;
        rom_memory[29724] = 3'b111;
        rom_memory[29725] = 3'b111;
        rom_memory[29726] = 3'b111;
        rom_memory[29727] = 3'b111;
        rom_memory[29728] = 3'b111;
        rom_memory[29729] = 3'b111;
        rom_memory[29730] = 3'b111;
        rom_memory[29731] = 3'b111;
        rom_memory[29732] = 3'b111;
        rom_memory[29733] = 3'b111;
        rom_memory[29734] = 3'b111;
        rom_memory[29735] = 3'b111;
        rom_memory[29736] = 3'b111;
        rom_memory[29737] = 3'b111;
        rom_memory[29738] = 3'b111;
        rom_memory[29739] = 3'b111;
        rom_memory[29740] = 3'b111;
        rom_memory[29741] = 3'b111;
        rom_memory[29742] = 3'b111;
        rom_memory[29743] = 3'b111;
        rom_memory[29744] = 3'b111;
        rom_memory[29745] = 3'b111;
        rom_memory[29746] = 3'b111;
        rom_memory[29747] = 3'b111;
        rom_memory[29748] = 3'b111;
        rom_memory[29749] = 3'b111;
        rom_memory[29750] = 3'b111;
        rom_memory[29751] = 3'b111;
        rom_memory[29752] = 3'b111;
        rom_memory[29753] = 3'b111;
        rom_memory[29754] = 3'b111;
        rom_memory[29755] = 3'b111;
        rom_memory[29756] = 3'b111;
        rom_memory[29757] = 3'b111;
        rom_memory[29758] = 3'b111;
        rom_memory[29759] = 3'b111;
        rom_memory[29760] = 3'b110;
        rom_memory[29761] = 3'b110;
        rom_memory[29762] = 3'b110;
        rom_memory[29763] = 3'b110;
        rom_memory[29764] = 3'b110;
        rom_memory[29765] = 3'b110;
        rom_memory[29766] = 3'b110;
        rom_memory[29767] = 3'b110;
        rom_memory[29768] = 3'b110;
        rom_memory[29769] = 3'b110;
        rom_memory[29770] = 3'b110;
        rom_memory[29771] = 3'b111;
        rom_memory[29772] = 3'b111;
        rom_memory[29773] = 3'b111;
        rom_memory[29774] = 3'b111;
        rom_memory[29775] = 3'b111;
        rom_memory[29776] = 3'b111;
        rom_memory[29777] = 3'b111;
        rom_memory[29778] = 3'b111;
        rom_memory[29779] = 3'b111;
        rom_memory[29780] = 3'b111;
        rom_memory[29781] = 3'b111;
        rom_memory[29782] = 3'b111;
        rom_memory[29783] = 3'b111;
        rom_memory[29784] = 3'b111;
        rom_memory[29785] = 3'b111;
        rom_memory[29786] = 3'b111;
        rom_memory[29787] = 3'b111;
        rom_memory[29788] = 3'b111;
        rom_memory[29789] = 3'b110;
        rom_memory[29790] = 3'b110;
        rom_memory[29791] = 3'b110;
        rom_memory[29792] = 3'b110;
        rom_memory[29793] = 3'b110;
        rom_memory[29794] = 3'b110;
        rom_memory[29795] = 3'b110;
        rom_memory[29796] = 3'b110;
        rom_memory[29797] = 3'b110;
        rom_memory[29798] = 3'b110;
        rom_memory[29799] = 3'b110;
        rom_memory[29800] = 3'b110;
        rom_memory[29801] = 3'b110;
        rom_memory[29802] = 3'b110;
        rom_memory[29803] = 3'b110;
        rom_memory[29804] = 3'b110;
        rom_memory[29805] = 3'b111;
        rom_memory[29806] = 3'b111;
        rom_memory[29807] = 3'b111;
        rom_memory[29808] = 3'b111;
        rom_memory[29809] = 3'b111;
        rom_memory[29810] = 3'b111;
        rom_memory[29811] = 3'b111;
        rom_memory[29812] = 3'b111;
        rom_memory[29813] = 3'b111;
        rom_memory[29814] = 3'b111;
        rom_memory[29815] = 3'b111;
        rom_memory[29816] = 3'b111;
        rom_memory[29817] = 3'b111;
        rom_memory[29818] = 3'b111;
        rom_memory[29819] = 3'b111;
        rom_memory[29820] = 3'b111;
        rom_memory[29821] = 3'b111;
        rom_memory[29822] = 3'b111;
        rom_memory[29823] = 3'b111;
        rom_memory[29824] = 3'b111;
        rom_memory[29825] = 3'b111;
        rom_memory[29826] = 3'b111;
        rom_memory[29827] = 3'b111;
        rom_memory[29828] = 3'b111;
        rom_memory[29829] = 3'b111;
        rom_memory[29830] = 3'b111;
        rom_memory[29831] = 3'b110;
        rom_memory[29832] = 3'b110;
        rom_memory[29833] = 3'b110;
        rom_memory[29834] = 3'b100;
        rom_memory[29835] = 3'b100;
        rom_memory[29836] = 3'b110;
        rom_memory[29837] = 3'b100;
        rom_memory[29838] = 3'b100;
        rom_memory[29839] = 3'b100;
        rom_memory[29840] = 3'b100;
        rom_memory[29841] = 3'b100;
        rom_memory[29842] = 3'b100;
        rom_memory[29843] = 3'b100;
        rom_memory[29844] = 3'b100;
        rom_memory[29845] = 3'b100;
        rom_memory[29846] = 3'b110;
        rom_memory[29847] = 3'b110;
        rom_memory[29848] = 3'b100;
        rom_memory[29849] = 3'b100;
        rom_memory[29850] = 3'b110;
        rom_memory[29851] = 3'b110;
        rom_memory[29852] = 3'b110;
        rom_memory[29853] = 3'b110;
        rom_memory[29854] = 3'b110;
        rom_memory[29855] = 3'b111;
        rom_memory[29856] = 3'b111;
        rom_memory[29857] = 3'b110;
        rom_memory[29858] = 3'b110;
        rom_memory[29859] = 3'b110;
        rom_memory[29860] = 3'b110;
        rom_memory[29861] = 3'b110;
        rom_memory[29862] = 3'b110;
        rom_memory[29863] = 3'b110;
        rom_memory[29864] = 3'b110;
        rom_memory[29865] = 3'b110;
        rom_memory[29866] = 3'b110;
        rom_memory[29867] = 3'b110;
        rom_memory[29868] = 3'b110;
        rom_memory[29869] = 3'b110;
        rom_memory[29870] = 3'b110;
        rom_memory[29871] = 3'b110;
        rom_memory[29872] = 3'b110;
        rom_memory[29873] = 3'b110;
        rom_memory[29874] = 3'b100;
        rom_memory[29875] = 3'b100;
        rom_memory[29876] = 3'b100;
        rom_memory[29877] = 3'b100;
        rom_memory[29878] = 3'b100;
        rom_memory[29879] = 3'b100;
        rom_memory[29880] = 3'b100;
        rom_memory[29881] = 3'b100;
        rom_memory[29882] = 3'b110;
        rom_memory[29883] = 3'b110;
        rom_memory[29884] = 3'b110;
        rom_memory[29885] = 3'b110;
        rom_memory[29886] = 3'b110;
        rom_memory[29887] = 3'b000;
        rom_memory[29888] = 3'b000;
        rom_memory[29889] = 3'b100;
        rom_memory[29890] = 3'b110;
        rom_memory[29891] = 3'b110;
        rom_memory[29892] = 3'b110;
        rom_memory[29893] = 3'b110;
        rom_memory[29894] = 3'b110;
        rom_memory[29895] = 3'b110;
        rom_memory[29896] = 3'b100;
        rom_memory[29897] = 3'b110;
        rom_memory[29898] = 3'b110;
        rom_memory[29899] = 3'b110;
        rom_memory[29900] = 3'b110;
        rom_memory[29901] = 3'b110;
        rom_memory[29902] = 3'b110;
        rom_memory[29903] = 3'b110;
        rom_memory[29904] = 3'b110;
        rom_memory[29905] = 3'b110;
        rom_memory[29906] = 3'b110;
        rom_memory[29907] = 3'b110;
        rom_memory[29908] = 3'b110;
        rom_memory[29909] = 3'b110;
        rom_memory[29910] = 3'b110;
        rom_memory[29911] = 3'b110;
        rom_memory[29912] = 3'b110;
        rom_memory[29913] = 3'b110;
        rom_memory[29914] = 3'b110;
        rom_memory[29915] = 3'b110;
        rom_memory[29916] = 3'b110;
        rom_memory[29917] = 3'b110;
        rom_memory[29918] = 3'b110;
        rom_memory[29919] = 3'b110;
        rom_memory[29920] = 3'b110;
        rom_memory[29921] = 3'b110;
        rom_memory[29922] = 3'b110;
        rom_memory[29923] = 3'b110;
        rom_memory[29924] = 3'b110;
        rom_memory[29925] = 3'b110;
        rom_memory[29926] = 3'b110;
        rom_memory[29927] = 3'b110;
        rom_memory[29928] = 3'b110;
        rom_memory[29929] = 3'b110;
        rom_memory[29930] = 3'b110;
        rom_memory[29931] = 3'b110;
        rom_memory[29932] = 3'b110;
        rom_memory[29933] = 3'b110;
        rom_memory[29934] = 3'b110;
        rom_memory[29935] = 3'b110;
        rom_memory[29936] = 3'b110;
        rom_memory[29937] = 3'b110;
        rom_memory[29938] = 3'b110;
        rom_memory[29939] = 3'b110;
        rom_memory[29940] = 3'b110;
        rom_memory[29941] = 3'b110;
        rom_memory[29942] = 3'b110;
        rom_memory[29943] = 3'b110;
        rom_memory[29944] = 3'b111;
        rom_memory[29945] = 3'b111;
        rom_memory[29946] = 3'b111;
        rom_memory[29947] = 3'b111;
        rom_memory[29948] = 3'b111;
        rom_memory[29949] = 3'b111;
        rom_memory[29950] = 3'b111;
        rom_memory[29951] = 3'b111;
        rom_memory[29952] = 3'b111;
        rom_memory[29953] = 3'b111;
        rom_memory[29954] = 3'b111;
        rom_memory[29955] = 3'b111;
        rom_memory[29956] = 3'b111;
        rom_memory[29957] = 3'b111;
        rom_memory[29958] = 3'b111;
        rom_memory[29959] = 3'b111;
        rom_memory[29960] = 3'b111;
        rom_memory[29961] = 3'b111;
        rom_memory[29962] = 3'b111;
        rom_memory[29963] = 3'b111;
        rom_memory[29964] = 3'b111;
        rom_memory[29965] = 3'b111;
        rom_memory[29966] = 3'b111;
        rom_memory[29967] = 3'b111;
        rom_memory[29968] = 3'b111;
        rom_memory[29969] = 3'b111;
        rom_memory[29970] = 3'b111;
        rom_memory[29971] = 3'b111;
        rom_memory[29972] = 3'b111;
        rom_memory[29973] = 3'b111;
        rom_memory[29974] = 3'b111;
        rom_memory[29975] = 3'b111;
        rom_memory[29976] = 3'b111;
        rom_memory[29977] = 3'b111;
        rom_memory[29978] = 3'b111;
        rom_memory[29979] = 3'b111;
        rom_memory[29980] = 3'b111;
        rom_memory[29981] = 3'b111;
        rom_memory[29982] = 3'b111;
        rom_memory[29983] = 3'b111;
        rom_memory[29984] = 3'b111;
        rom_memory[29985] = 3'b111;
        rom_memory[29986] = 3'b111;
        rom_memory[29987] = 3'b111;
        rom_memory[29988] = 3'b111;
        rom_memory[29989] = 3'b111;
        rom_memory[29990] = 3'b111;
        rom_memory[29991] = 3'b111;
        rom_memory[29992] = 3'b111;
        rom_memory[29993] = 3'b111;
        rom_memory[29994] = 3'b111;
        rom_memory[29995] = 3'b111;
        rom_memory[29996] = 3'b111;
        rom_memory[29997] = 3'b111;
        rom_memory[29998] = 3'b111;
        rom_memory[29999] = 3'b111;
        rom_memory[30000] = 3'b110;
        rom_memory[30001] = 3'b110;
        rom_memory[30002] = 3'b110;
        rom_memory[30003] = 3'b110;
        rom_memory[30004] = 3'b110;
        rom_memory[30005] = 3'b110;
        rom_memory[30006] = 3'b110;
        rom_memory[30007] = 3'b110;
        rom_memory[30008] = 3'b110;
        rom_memory[30009] = 3'b110;
        rom_memory[30010] = 3'b110;
        rom_memory[30011] = 3'b111;
        rom_memory[30012] = 3'b111;
        rom_memory[30013] = 3'b111;
        rom_memory[30014] = 3'b111;
        rom_memory[30015] = 3'b111;
        rom_memory[30016] = 3'b111;
        rom_memory[30017] = 3'b111;
        rom_memory[30018] = 3'b111;
        rom_memory[30019] = 3'b111;
        rom_memory[30020] = 3'b111;
        rom_memory[30021] = 3'b111;
        rom_memory[30022] = 3'b111;
        rom_memory[30023] = 3'b111;
        rom_memory[30024] = 3'b111;
        rom_memory[30025] = 3'b111;
        rom_memory[30026] = 3'b111;
        rom_memory[30027] = 3'b111;
        rom_memory[30028] = 3'b111;
        rom_memory[30029] = 3'b110;
        rom_memory[30030] = 3'b110;
        rom_memory[30031] = 3'b110;
        rom_memory[30032] = 3'b110;
        rom_memory[30033] = 3'b111;
        rom_memory[30034] = 3'b111;
        rom_memory[30035] = 3'b111;
        rom_memory[30036] = 3'b110;
        rom_memory[30037] = 3'b110;
        rom_memory[30038] = 3'b110;
        rom_memory[30039] = 3'b110;
        rom_memory[30040] = 3'b110;
        rom_memory[30041] = 3'b110;
        rom_memory[30042] = 3'b110;
        rom_memory[30043] = 3'b110;
        rom_memory[30044] = 3'b110;
        rom_memory[30045] = 3'b111;
        rom_memory[30046] = 3'b111;
        rom_memory[30047] = 3'b111;
        rom_memory[30048] = 3'b111;
        rom_memory[30049] = 3'b111;
        rom_memory[30050] = 3'b111;
        rom_memory[30051] = 3'b111;
        rom_memory[30052] = 3'b111;
        rom_memory[30053] = 3'b111;
        rom_memory[30054] = 3'b111;
        rom_memory[30055] = 3'b111;
        rom_memory[30056] = 3'b111;
        rom_memory[30057] = 3'b111;
        rom_memory[30058] = 3'b111;
        rom_memory[30059] = 3'b111;
        rom_memory[30060] = 3'b111;
        rom_memory[30061] = 3'b111;
        rom_memory[30062] = 3'b111;
        rom_memory[30063] = 3'b111;
        rom_memory[30064] = 3'b111;
        rom_memory[30065] = 3'b111;
        rom_memory[30066] = 3'b111;
        rom_memory[30067] = 3'b111;
        rom_memory[30068] = 3'b111;
        rom_memory[30069] = 3'b111;
        rom_memory[30070] = 3'b111;
        rom_memory[30071] = 3'b111;
        rom_memory[30072] = 3'b111;
        rom_memory[30073] = 3'b111;
        rom_memory[30074] = 3'b110;
        rom_memory[30075] = 3'b110;
        rom_memory[30076] = 3'b110;
        rom_memory[30077] = 3'b110;
        rom_memory[30078] = 3'b100;
        rom_memory[30079] = 3'b100;
        rom_memory[30080] = 3'b100;
        rom_memory[30081] = 3'b110;
        rom_memory[30082] = 3'b100;
        rom_memory[30083] = 3'b100;
        rom_memory[30084] = 3'b100;
        rom_memory[30085] = 3'b100;
        rom_memory[30086] = 3'b100;
        rom_memory[30087] = 3'b100;
        rom_memory[30088] = 3'b100;
        rom_memory[30089] = 3'b100;
        rom_memory[30090] = 3'b110;
        rom_memory[30091] = 3'b111;
        rom_memory[30092] = 3'b111;
        rom_memory[30093] = 3'b110;
        rom_memory[30094] = 3'b110;
        rom_memory[30095] = 3'b111;
        rom_memory[30096] = 3'b111;
        rom_memory[30097] = 3'b110;
        rom_memory[30098] = 3'b110;
        rom_memory[30099] = 3'b100;
        rom_memory[30100] = 3'b110;
        rom_memory[30101] = 3'b110;
        rom_memory[30102] = 3'b110;
        rom_memory[30103] = 3'b110;
        rom_memory[30104] = 3'b110;
        rom_memory[30105] = 3'b110;
        rom_memory[30106] = 3'b110;
        rom_memory[30107] = 3'b110;
        rom_memory[30108] = 3'b110;
        rom_memory[30109] = 3'b110;
        rom_memory[30110] = 3'b110;
        rom_memory[30111] = 3'b110;
        rom_memory[30112] = 3'b110;
        rom_memory[30113] = 3'b110;
        rom_memory[30114] = 3'b110;
        rom_memory[30115] = 3'b100;
        rom_memory[30116] = 3'b100;
        rom_memory[30117] = 3'b100;
        rom_memory[30118] = 3'b100;
        rom_memory[30119] = 3'b100;
        rom_memory[30120] = 3'b100;
        rom_memory[30121] = 3'b100;
        rom_memory[30122] = 3'b100;
        rom_memory[30123] = 3'b100;
        rom_memory[30124] = 3'b110;
        rom_memory[30125] = 3'b110;
        rom_memory[30126] = 3'b110;
        rom_memory[30127] = 3'b100;
        rom_memory[30128] = 3'b000;
        rom_memory[30129] = 3'b000;
        rom_memory[30130] = 3'b100;
        rom_memory[30131] = 3'b110;
        rom_memory[30132] = 3'b110;
        rom_memory[30133] = 3'b110;
        rom_memory[30134] = 3'b110;
        rom_memory[30135] = 3'b100;
        rom_memory[30136] = 3'b100;
        rom_memory[30137] = 3'b100;
        rom_memory[30138] = 3'b110;
        rom_memory[30139] = 3'b111;
        rom_memory[30140] = 3'b110;
        rom_memory[30141] = 3'b110;
        rom_memory[30142] = 3'b110;
        rom_memory[30143] = 3'b110;
        rom_memory[30144] = 3'b110;
        rom_memory[30145] = 3'b110;
        rom_memory[30146] = 3'b110;
        rom_memory[30147] = 3'b110;
        rom_memory[30148] = 3'b110;
        rom_memory[30149] = 3'b110;
        rom_memory[30150] = 3'b110;
        rom_memory[30151] = 3'b110;
        rom_memory[30152] = 3'b110;
        rom_memory[30153] = 3'b110;
        rom_memory[30154] = 3'b110;
        rom_memory[30155] = 3'b110;
        rom_memory[30156] = 3'b110;
        rom_memory[30157] = 3'b110;
        rom_memory[30158] = 3'b110;
        rom_memory[30159] = 3'b110;
        rom_memory[30160] = 3'b110;
        rom_memory[30161] = 3'b110;
        rom_memory[30162] = 3'b110;
        rom_memory[30163] = 3'b110;
        rom_memory[30164] = 3'b110;
        rom_memory[30165] = 3'b110;
        rom_memory[30166] = 3'b110;
        rom_memory[30167] = 3'b110;
        rom_memory[30168] = 3'b110;
        rom_memory[30169] = 3'b110;
        rom_memory[30170] = 3'b110;
        rom_memory[30171] = 3'b110;
        rom_memory[30172] = 3'b110;
        rom_memory[30173] = 3'b110;
        rom_memory[30174] = 3'b110;
        rom_memory[30175] = 3'b110;
        rom_memory[30176] = 3'b110;
        rom_memory[30177] = 3'b110;
        rom_memory[30178] = 3'b110;
        rom_memory[30179] = 3'b110;
        rom_memory[30180] = 3'b110;
        rom_memory[30181] = 3'b110;
        rom_memory[30182] = 3'b110;
        rom_memory[30183] = 3'b110;
        rom_memory[30184] = 3'b111;
        rom_memory[30185] = 3'b111;
        rom_memory[30186] = 3'b111;
        rom_memory[30187] = 3'b111;
        rom_memory[30188] = 3'b111;
        rom_memory[30189] = 3'b111;
        rom_memory[30190] = 3'b111;
        rom_memory[30191] = 3'b111;
        rom_memory[30192] = 3'b111;
        rom_memory[30193] = 3'b111;
        rom_memory[30194] = 3'b111;
        rom_memory[30195] = 3'b111;
        rom_memory[30196] = 3'b111;
        rom_memory[30197] = 3'b111;
        rom_memory[30198] = 3'b111;
        rom_memory[30199] = 3'b111;
        rom_memory[30200] = 3'b111;
        rom_memory[30201] = 3'b111;
        rom_memory[30202] = 3'b111;
        rom_memory[30203] = 3'b111;
        rom_memory[30204] = 3'b111;
        rom_memory[30205] = 3'b111;
        rom_memory[30206] = 3'b111;
        rom_memory[30207] = 3'b111;
        rom_memory[30208] = 3'b111;
        rom_memory[30209] = 3'b111;
        rom_memory[30210] = 3'b111;
        rom_memory[30211] = 3'b111;
        rom_memory[30212] = 3'b111;
        rom_memory[30213] = 3'b111;
        rom_memory[30214] = 3'b111;
        rom_memory[30215] = 3'b111;
        rom_memory[30216] = 3'b111;
        rom_memory[30217] = 3'b111;
        rom_memory[30218] = 3'b111;
        rom_memory[30219] = 3'b111;
        rom_memory[30220] = 3'b111;
        rom_memory[30221] = 3'b111;
        rom_memory[30222] = 3'b111;
        rom_memory[30223] = 3'b111;
        rom_memory[30224] = 3'b111;
        rom_memory[30225] = 3'b111;
        rom_memory[30226] = 3'b111;
        rom_memory[30227] = 3'b111;
        rom_memory[30228] = 3'b111;
        rom_memory[30229] = 3'b111;
        rom_memory[30230] = 3'b111;
        rom_memory[30231] = 3'b111;
        rom_memory[30232] = 3'b111;
        rom_memory[30233] = 3'b111;
        rom_memory[30234] = 3'b111;
        rom_memory[30235] = 3'b111;
        rom_memory[30236] = 3'b111;
        rom_memory[30237] = 3'b111;
        rom_memory[30238] = 3'b111;
        rom_memory[30239] = 3'b111;
        rom_memory[30240] = 3'b110;
        rom_memory[30241] = 3'b110;
        rom_memory[30242] = 3'b110;
        rom_memory[30243] = 3'b110;
        rom_memory[30244] = 3'b110;
        rom_memory[30245] = 3'b110;
        rom_memory[30246] = 3'b110;
        rom_memory[30247] = 3'b110;
        rom_memory[30248] = 3'b110;
        rom_memory[30249] = 3'b110;
        rom_memory[30250] = 3'b110;
        rom_memory[30251] = 3'b111;
        rom_memory[30252] = 3'b111;
        rom_memory[30253] = 3'b111;
        rom_memory[30254] = 3'b111;
        rom_memory[30255] = 3'b111;
        rom_memory[30256] = 3'b111;
        rom_memory[30257] = 3'b111;
        rom_memory[30258] = 3'b111;
        rom_memory[30259] = 3'b111;
        rom_memory[30260] = 3'b111;
        rom_memory[30261] = 3'b111;
        rom_memory[30262] = 3'b111;
        rom_memory[30263] = 3'b111;
        rom_memory[30264] = 3'b111;
        rom_memory[30265] = 3'b111;
        rom_memory[30266] = 3'b111;
        rom_memory[30267] = 3'b111;
        rom_memory[30268] = 3'b111;
        rom_memory[30269] = 3'b110;
        rom_memory[30270] = 3'b110;
        rom_memory[30271] = 3'b110;
        rom_memory[30272] = 3'b111;
        rom_memory[30273] = 3'b111;
        rom_memory[30274] = 3'b111;
        rom_memory[30275] = 3'b111;
        rom_memory[30276] = 3'b110;
        rom_memory[30277] = 3'b110;
        rom_memory[30278] = 3'b110;
        rom_memory[30279] = 3'b110;
        rom_memory[30280] = 3'b110;
        rom_memory[30281] = 3'b110;
        rom_memory[30282] = 3'b110;
        rom_memory[30283] = 3'b110;
        rom_memory[30284] = 3'b110;
        rom_memory[30285] = 3'b110;
        rom_memory[30286] = 3'b110;
        rom_memory[30287] = 3'b110;
        rom_memory[30288] = 3'b110;
        rom_memory[30289] = 3'b111;
        rom_memory[30290] = 3'b111;
        rom_memory[30291] = 3'b111;
        rom_memory[30292] = 3'b111;
        rom_memory[30293] = 3'b111;
        rom_memory[30294] = 3'b111;
        rom_memory[30295] = 3'b111;
        rom_memory[30296] = 3'b111;
        rom_memory[30297] = 3'b111;
        rom_memory[30298] = 3'b111;
        rom_memory[30299] = 3'b111;
        rom_memory[30300] = 3'b111;
        rom_memory[30301] = 3'b111;
        rom_memory[30302] = 3'b111;
        rom_memory[30303] = 3'b111;
        rom_memory[30304] = 3'b111;
        rom_memory[30305] = 3'b111;
        rom_memory[30306] = 3'b111;
        rom_memory[30307] = 3'b111;
        rom_memory[30308] = 3'b111;
        rom_memory[30309] = 3'b111;
        rom_memory[30310] = 3'b111;
        rom_memory[30311] = 3'b111;
        rom_memory[30312] = 3'b111;
        rom_memory[30313] = 3'b111;
        rom_memory[30314] = 3'b111;
        rom_memory[30315] = 3'b110;
        rom_memory[30316] = 3'b110;
        rom_memory[30317] = 3'b110;
        rom_memory[30318] = 3'b110;
        rom_memory[30319] = 3'b110;
        rom_memory[30320] = 3'b110;
        rom_memory[30321] = 3'b111;
        rom_memory[30322] = 3'b110;
        rom_memory[30323] = 3'b100;
        rom_memory[30324] = 3'b000;
        rom_memory[30325] = 3'b000;
        rom_memory[30326] = 3'b000;
        rom_memory[30327] = 3'b100;
        rom_memory[30328] = 3'b100;
        rom_memory[30329] = 3'b100;
        rom_memory[30330] = 3'b110;
        rom_memory[30331] = 3'b110;
        rom_memory[30332] = 3'b111;
        rom_memory[30333] = 3'b110;
        rom_memory[30334] = 3'b111;
        rom_memory[30335] = 3'b111;
        rom_memory[30336] = 3'b110;
        rom_memory[30337] = 3'b110;
        rom_memory[30338] = 3'b110;
        rom_memory[30339] = 3'b100;
        rom_memory[30340] = 3'b100;
        rom_memory[30341] = 3'b000;
        rom_memory[30342] = 3'b100;
        rom_memory[30343] = 3'b110;
        rom_memory[30344] = 3'b110;
        rom_memory[30345] = 3'b110;
        rom_memory[30346] = 3'b110;
        rom_memory[30347] = 3'b110;
        rom_memory[30348] = 3'b110;
        rom_memory[30349] = 3'b110;
        rom_memory[30350] = 3'b111;
        rom_memory[30351] = 3'b110;
        rom_memory[30352] = 3'b110;
        rom_memory[30353] = 3'b110;
        rom_memory[30354] = 3'b110;
        rom_memory[30355] = 3'b110;
        rom_memory[30356] = 3'b110;
        rom_memory[30357] = 3'b110;
        rom_memory[30358] = 3'b110;
        rom_memory[30359] = 3'b100;
        rom_memory[30360] = 3'b100;
        rom_memory[30361] = 3'b100;
        rom_memory[30362] = 3'b100;
        rom_memory[30363] = 3'b100;
        rom_memory[30364] = 3'b100;
        rom_memory[30365] = 3'b100;
        rom_memory[30366] = 3'b100;
        rom_memory[30367] = 3'b100;
        rom_memory[30368] = 3'b100;
        rom_memory[30369] = 3'b000;
        rom_memory[30370] = 3'b000;
        rom_memory[30371] = 3'b100;
        rom_memory[30372] = 3'b110;
        rom_memory[30373] = 3'b110;
        rom_memory[30374] = 3'b110;
        rom_memory[30375] = 3'b110;
        rom_memory[30376] = 3'b100;
        rom_memory[30377] = 3'b110;
        rom_memory[30378] = 3'b100;
        rom_memory[30379] = 3'b110;
        rom_memory[30380] = 3'b111;
        rom_memory[30381] = 3'b110;
        rom_memory[30382] = 3'b110;
        rom_memory[30383] = 3'b110;
        rom_memory[30384] = 3'b110;
        rom_memory[30385] = 3'b110;
        rom_memory[30386] = 3'b110;
        rom_memory[30387] = 3'b110;
        rom_memory[30388] = 3'b110;
        rom_memory[30389] = 3'b110;
        rom_memory[30390] = 3'b110;
        rom_memory[30391] = 3'b110;
        rom_memory[30392] = 3'b110;
        rom_memory[30393] = 3'b110;
        rom_memory[30394] = 3'b110;
        rom_memory[30395] = 3'b110;
        rom_memory[30396] = 3'b110;
        rom_memory[30397] = 3'b110;
        rom_memory[30398] = 3'b110;
        rom_memory[30399] = 3'b110;
        rom_memory[30400] = 3'b110;
        rom_memory[30401] = 3'b110;
        rom_memory[30402] = 3'b110;
        rom_memory[30403] = 3'b110;
        rom_memory[30404] = 3'b110;
        rom_memory[30405] = 3'b110;
        rom_memory[30406] = 3'b110;
        rom_memory[30407] = 3'b110;
        rom_memory[30408] = 3'b110;
        rom_memory[30409] = 3'b110;
        rom_memory[30410] = 3'b110;
        rom_memory[30411] = 3'b110;
        rom_memory[30412] = 3'b110;
        rom_memory[30413] = 3'b110;
        rom_memory[30414] = 3'b110;
        rom_memory[30415] = 3'b110;
        rom_memory[30416] = 3'b110;
        rom_memory[30417] = 3'b110;
        rom_memory[30418] = 3'b110;
        rom_memory[30419] = 3'b110;
        rom_memory[30420] = 3'b110;
        rom_memory[30421] = 3'b110;
        rom_memory[30422] = 3'b110;
        rom_memory[30423] = 3'b110;
        rom_memory[30424] = 3'b111;
        rom_memory[30425] = 3'b111;
        rom_memory[30426] = 3'b111;
        rom_memory[30427] = 3'b111;
        rom_memory[30428] = 3'b111;
        rom_memory[30429] = 3'b111;
        rom_memory[30430] = 3'b111;
        rom_memory[30431] = 3'b111;
        rom_memory[30432] = 3'b111;
        rom_memory[30433] = 3'b111;
        rom_memory[30434] = 3'b111;
        rom_memory[30435] = 3'b111;
        rom_memory[30436] = 3'b111;
        rom_memory[30437] = 3'b111;
        rom_memory[30438] = 3'b111;
        rom_memory[30439] = 3'b111;
        rom_memory[30440] = 3'b111;
        rom_memory[30441] = 3'b111;
        rom_memory[30442] = 3'b111;
        rom_memory[30443] = 3'b111;
        rom_memory[30444] = 3'b111;
        rom_memory[30445] = 3'b111;
        rom_memory[30446] = 3'b111;
        rom_memory[30447] = 3'b111;
        rom_memory[30448] = 3'b111;
        rom_memory[30449] = 3'b111;
        rom_memory[30450] = 3'b111;
        rom_memory[30451] = 3'b111;
        rom_memory[30452] = 3'b111;
        rom_memory[30453] = 3'b111;
        rom_memory[30454] = 3'b111;
        rom_memory[30455] = 3'b111;
        rom_memory[30456] = 3'b111;
        rom_memory[30457] = 3'b111;
        rom_memory[30458] = 3'b111;
        rom_memory[30459] = 3'b111;
        rom_memory[30460] = 3'b111;
        rom_memory[30461] = 3'b111;
        rom_memory[30462] = 3'b111;
        rom_memory[30463] = 3'b111;
        rom_memory[30464] = 3'b111;
        rom_memory[30465] = 3'b111;
        rom_memory[30466] = 3'b111;
        rom_memory[30467] = 3'b111;
        rom_memory[30468] = 3'b111;
        rom_memory[30469] = 3'b111;
        rom_memory[30470] = 3'b111;
        rom_memory[30471] = 3'b111;
        rom_memory[30472] = 3'b111;
        rom_memory[30473] = 3'b111;
        rom_memory[30474] = 3'b111;
        rom_memory[30475] = 3'b111;
        rom_memory[30476] = 3'b111;
        rom_memory[30477] = 3'b111;
        rom_memory[30478] = 3'b111;
        rom_memory[30479] = 3'b111;
        rom_memory[30480] = 3'b110;
        rom_memory[30481] = 3'b110;
        rom_memory[30482] = 3'b110;
        rom_memory[30483] = 3'b110;
        rom_memory[30484] = 3'b110;
        rom_memory[30485] = 3'b110;
        rom_memory[30486] = 3'b110;
        rom_memory[30487] = 3'b110;
        rom_memory[30488] = 3'b110;
        rom_memory[30489] = 3'b110;
        rom_memory[30490] = 3'b110;
        rom_memory[30491] = 3'b110;
        rom_memory[30492] = 3'b111;
        rom_memory[30493] = 3'b111;
        rom_memory[30494] = 3'b111;
        rom_memory[30495] = 3'b111;
        rom_memory[30496] = 3'b111;
        rom_memory[30497] = 3'b111;
        rom_memory[30498] = 3'b111;
        rom_memory[30499] = 3'b111;
        rom_memory[30500] = 3'b111;
        rom_memory[30501] = 3'b111;
        rom_memory[30502] = 3'b111;
        rom_memory[30503] = 3'b111;
        rom_memory[30504] = 3'b111;
        rom_memory[30505] = 3'b111;
        rom_memory[30506] = 3'b111;
        rom_memory[30507] = 3'b111;
        rom_memory[30508] = 3'b111;
        rom_memory[30509] = 3'b111;
        rom_memory[30510] = 3'b111;
        rom_memory[30511] = 3'b111;
        rom_memory[30512] = 3'b111;
        rom_memory[30513] = 3'b111;
        rom_memory[30514] = 3'b111;
        rom_memory[30515] = 3'b111;
        rom_memory[30516] = 3'b110;
        rom_memory[30517] = 3'b110;
        rom_memory[30518] = 3'b110;
        rom_memory[30519] = 3'b110;
        rom_memory[30520] = 3'b110;
        rom_memory[30521] = 3'b110;
        rom_memory[30522] = 3'b110;
        rom_memory[30523] = 3'b110;
        rom_memory[30524] = 3'b110;
        rom_memory[30525] = 3'b110;
        rom_memory[30526] = 3'b111;
        rom_memory[30527] = 3'b111;
        rom_memory[30528] = 3'b111;
        rom_memory[30529] = 3'b111;
        rom_memory[30530] = 3'b111;
        rom_memory[30531] = 3'b111;
        rom_memory[30532] = 3'b111;
        rom_memory[30533] = 3'b111;
        rom_memory[30534] = 3'b111;
        rom_memory[30535] = 3'b111;
        rom_memory[30536] = 3'b111;
        rom_memory[30537] = 3'b111;
        rom_memory[30538] = 3'b111;
        rom_memory[30539] = 3'b111;
        rom_memory[30540] = 3'b111;
        rom_memory[30541] = 3'b111;
        rom_memory[30542] = 3'b111;
        rom_memory[30543] = 3'b111;
        rom_memory[30544] = 3'b111;
        rom_memory[30545] = 3'b111;
        rom_memory[30546] = 3'b111;
        rom_memory[30547] = 3'b111;
        rom_memory[30548] = 3'b110;
        rom_memory[30549] = 3'b110;
        rom_memory[30550] = 3'b110;
        rom_memory[30551] = 3'b110;
        rom_memory[30552] = 3'b110;
        rom_memory[30553] = 3'b110;
        rom_memory[30554] = 3'b110;
        rom_memory[30555] = 3'b111;
        rom_memory[30556] = 3'b111;
        rom_memory[30557] = 3'b110;
        rom_memory[30558] = 3'b110;
        rom_memory[30559] = 3'b110;
        rom_memory[30560] = 3'b110;
        rom_memory[30561] = 3'b111;
        rom_memory[30562] = 3'b111;
        rom_memory[30563] = 3'b000;
        rom_memory[30564] = 3'b000;
        rom_memory[30565] = 3'b100;
        rom_memory[30566] = 3'b000;
        rom_memory[30567] = 3'b000;
        rom_memory[30568] = 3'b100;
        rom_memory[30569] = 3'b100;
        rom_memory[30570] = 3'b110;
        rom_memory[30571] = 3'b100;
        rom_memory[30572] = 3'b111;
        rom_memory[30573] = 3'b111;
        rom_memory[30574] = 3'b111;
        rom_memory[30575] = 3'b110;
        rom_memory[30576] = 3'b110;
        rom_memory[30577] = 3'b111;
        rom_memory[30578] = 3'b110;
        rom_memory[30579] = 3'b110;
        rom_memory[30580] = 3'b110;
        rom_memory[30581] = 3'b000;
        rom_memory[30582] = 3'b110;
        rom_memory[30583] = 3'b110;
        rom_memory[30584] = 3'b110;
        rom_memory[30585] = 3'b110;
        rom_memory[30586] = 3'b110;
        rom_memory[30587] = 3'b110;
        rom_memory[30588] = 3'b110;
        rom_memory[30589] = 3'b110;
        rom_memory[30590] = 3'b110;
        rom_memory[30591] = 3'b110;
        rom_memory[30592] = 3'b110;
        rom_memory[30593] = 3'b110;
        rom_memory[30594] = 3'b110;
        rom_memory[30595] = 3'b110;
        rom_memory[30596] = 3'b110;
        rom_memory[30597] = 3'b110;
        rom_memory[30598] = 3'b110;
        rom_memory[30599] = 3'b110;
        rom_memory[30600] = 3'b110;
        rom_memory[30601] = 3'b110;
        rom_memory[30602] = 3'b100;
        rom_memory[30603] = 3'b100;
        rom_memory[30604] = 3'b100;
        rom_memory[30605] = 3'b100;
        rom_memory[30606] = 3'b100;
        rom_memory[30607] = 3'b100;
        rom_memory[30608] = 3'b100;
        rom_memory[30609] = 3'b000;
        rom_memory[30610] = 3'b000;
        rom_memory[30611] = 3'b000;
        rom_memory[30612] = 3'b100;
        rom_memory[30613] = 3'b110;
        rom_memory[30614] = 3'b110;
        rom_memory[30615] = 3'b110;
        rom_memory[30616] = 3'b110;
        rom_memory[30617] = 3'b100;
        rom_memory[30618] = 3'b110;
        rom_memory[30619] = 3'b100;
        rom_memory[30620] = 3'b110;
        rom_memory[30621] = 3'b111;
        rom_memory[30622] = 3'b110;
        rom_memory[30623] = 3'b110;
        rom_memory[30624] = 3'b110;
        rom_memory[30625] = 3'b110;
        rom_memory[30626] = 3'b110;
        rom_memory[30627] = 3'b110;
        rom_memory[30628] = 3'b110;
        rom_memory[30629] = 3'b110;
        rom_memory[30630] = 3'b110;
        rom_memory[30631] = 3'b110;
        rom_memory[30632] = 3'b110;
        rom_memory[30633] = 3'b110;
        rom_memory[30634] = 3'b110;
        rom_memory[30635] = 3'b110;
        rom_memory[30636] = 3'b110;
        rom_memory[30637] = 3'b110;
        rom_memory[30638] = 3'b110;
        rom_memory[30639] = 3'b110;
        rom_memory[30640] = 3'b110;
        rom_memory[30641] = 3'b110;
        rom_memory[30642] = 3'b110;
        rom_memory[30643] = 3'b110;
        rom_memory[30644] = 3'b110;
        rom_memory[30645] = 3'b110;
        rom_memory[30646] = 3'b110;
        rom_memory[30647] = 3'b110;
        rom_memory[30648] = 3'b110;
        rom_memory[30649] = 3'b110;
        rom_memory[30650] = 3'b110;
        rom_memory[30651] = 3'b110;
        rom_memory[30652] = 3'b110;
        rom_memory[30653] = 3'b110;
        rom_memory[30654] = 3'b110;
        rom_memory[30655] = 3'b110;
        rom_memory[30656] = 3'b110;
        rom_memory[30657] = 3'b110;
        rom_memory[30658] = 3'b110;
        rom_memory[30659] = 3'b110;
        rom_memory[30660] = 3'b110;
        rom_memory[30661] = 3'b110;
        rom_memory[30662] = 3'b110;
        rom_memory[30663] = 3'b110;
        rom_memory[30664] = 3'b111;
        rom_memory[30665] = 3'b111;
        rom_memory[30666] = 3'b111;
        rom_memory[30667] = 3'b111;
        rom_memory[30668] = 3'b111;
        rom_memory[30669] = 3'b111;
        rom_memory[30670] = 3'b111;
        rom_memory[30671] = 3'b111;
        rom_memory[30672] = 3'b111;
        rom_memory[30673] = 3'b111;
        rom_memory[30674] = 3'b111;
        rom_memory[30675] = 3'b111;
        rom_memory[30676] = 3'b111;
        rom_memory[30677] = 3'b111;
        rom_memory[30678] = 3'b111;
        rom_memory[30679] = 3'b111;
        rom_memory[30680] = 3'b111;
        rom_memory[30681] = 3'b111;
        rom_memory[30682] = 3'b111;
        rom_memory[30683] = 3'b111;
        rom_memory[30684] = 3'b111;
        rom_memory[30685] = 3'b111;
        rom_memory[30686] = 3'b111;
        rom_memory[30687] = 3'b111;
        rom_memory[30688] = 3'b111;
        rom_memory[30689] = 3'b111;
        rom_memory[30690] = 3'b111;
        rom_memory[30691] = 3'b111;
        rom_memory[30692] = 3'b111;
        rom_memory[30693] = 3'b111;
        rom_memory[30694] = 3'b111;
        rom_memory[30695] = 3'b111;
        rom_memory[30696] = 3'b111;
        rom_memory[30697] = 3'b111;
        rom_memory[30698] = 3'b111;
        rom_memory[30699] = 3'b111;
        rom_memory[30700] = 3'b111;
        rom_memory[30701] = 3'b111;
        rom_memory[30702] = 3'b111;
        rom_memory[30703] = 3'b111;
        rom_memory[30704] = 3'b111;
        rom_memory[30705] = 3'b111;
        rom_memory[30706] = 3'b111;
        rom_memory[30707] = 3'b111;
        rom_memory[30708] = 3'b111;
        rom_memory[30709] = 3'b111;
        rom_memory[30710] = 3'b111;
        rom_memory[30711] = 3'b111;
        rom_memory[30712] = 3'b111;
        rom_memory[30713] = 3'b111;
        rom_memory[30714] = 3'b111;
        rom_memory[30715] = 3'b111;
        rom_memory[30716] = 3'b111;
        rom_memory[30717] = 3'b111;
        rom_memory[30718] = 3'b111;
        rom_memory[30719] = 3'b111;
        rom_memory[30720] = 3'b110;
        rom_memory[30721] = 3'b110;
        rom_memory[30722] = 3'b110;
        rom_memory[30723] = 3'b110;
        rom_memory[30724] = 3'b110;
        rom_memory[30725] = 3'b110;
        rom_memory[30726] = 3'b110;
        rom_memory[30727] = 3'b110;
        rom_memory[30728] = 3'b110;
        rom_memory[30729] = 3'b110;
        rom_memory[30730] = 3'b110;
        rom_memory[30731] = 3'b110;
        rom_memory[30732] = 3'b111;
        rom_memory[30733] = 3'b111;
        rom_memory[30734] = 3'b111;
        rom_memory[30735] = 3'b111;
        rom_memory[30736] = 3'b111;
        rom_memory[30737] = 3'b111;
        rom_memory[30738] = 3'b111;
        rom_memory[30739] = 3'b111;
        rom_memory[30740] = 3'b111;
        rom_memory[30741] = 3'b111;
        rom_memory[30742] = 3'b111;
        rom_memory[30743] = 3'b111;
        rom_memory[30744] = 3'b111;
        rom_memory[30745] = 3'b111;
        rom_memory[30746] = 3'b111;
        rom_memory[30747] = 3'b111;
        rom_memory[30748] = 3'b111;
        rom_memory[30749] = 3'b111;
        rom_memory[30750] = 3'b111;
        rom_memory[30751] = 3'b111;
        rom_memory[30752] = 3'b111;
        rom_memory[30753] = 3'b111;
        rom_memory[30754] = 3'b111;
        rom_memory[30755] = 3'b111;
        rom_memory[30756] = 3'b110;
        rom_memory[30757] = 3'b110;
        rom_memory[30758] = 3'b110;
        rom_memory[30759] = 3'b111;
        rom_memory[30760] = 3'b111;
        rom_memory[30761] = 3'b110;
        rom_memory[30762] = 3'b110;
        rom_memory[30763] = 3'b110;
        rom_memory[30764] = 3'b110;
        rom_memory[30765] = 3'b110;
        rom_memory[30766] = 3'b111;
        rom_memory[30767] = 3'b111;
        rom_memory[30768] = 3'b111;
        rom_memory[30769] = 3'b111;
        rom_memory[30770] = 3'b111;
        rom_memory[30771] = 3'b111;
        rom_memory[30772] = 3'b111;
        rom_memory[30773] = 3'b111;
        rom_memory[30774] = 3'b111;
        rom_memory[30775] = 3'b111;
        rom_memory[30776] = 3'b111;
        rom_memory[30777] = 3'b111;
        rom_memory[30778] = 3'b111;
        rom_memory[30779] = 3'b111;
        rom_memory[30780] = 3'b111;
        rom_memory[30781] = 3'b111;
        rom_memory[30782] = 3'b111;
        rom_memory[30783] = 3'b111;
        rom_memory[30784] = 3'b111;
        rom_memory[30785] = 3'b111;
        rom_memory[30786] = 3'b110;
        rom_memory[30787] = 3'b110;
        rom_memory[30788] = 3'b110;
        rom_memory[30789] = 3'b110;
        rom_memory[30790] = 3'b110;
        rom_memory[30791] = 3'b110;
        rom_memory[30792] = 3'b110;
        rom_memory[30793] = 3'b110;
        rom_memory[30794] = 3'b110;
        rom_memory[30795] = 3'b110;
        rom_memory[30796] = 3'b110;
        rom_memory[30797] = 3'b110;
        rom_memory[30798] = 3'b110;
        rom_memory[30799] = 3'b110;
        rom_memory[30800] = 3'b110;
        rom_memory[30801] = 3'b111;
        rom_memory[30802] = 3'b111;
        rom_memory[30803] = 3'b110;
        rom_memory[30804] = 3'b000;
        rom_memory[30805] = 3'b100;
        rom_memory[30806] = 3'b000;
        rom_memory[30807] = 3'b000;
        rom_memory[30808] = 3'b000;
        rom_memory[30809] = 3'b000;
        rom_memory[30810] = 3'b110;
        rom_memory[30811] = 3'b110;
        rom_memory[30812] = 3'b100;
        rom_memory[30813] = 3'b110;
        rom_memory[30814] = 3'b110;
        rom_memory[30815] = 3'b110;
        rom_memory[30816] = 3'b111;
        rom_memory[30817] = 3'b110;
        rom_memory[30818] = 3'b100;
        rom_memory[30819] = 3'b100;
        rom_memory[30820] = 3'b110;
        rom_memory[30821] = 3'b110;
        rom_memory[30822] = 3'b110;
        rom_memory[30823] = 3'b110;
        rom_memory[30824] = 3'b110;
        rom_memory[30825] = 3'b110;
        rom_memory[30826] = 3'b110;
        rom_memory[30827] = 3'b110;
        rom_memory[30828] = 3'b110;
        rom_memory[30829] = 3'b110;
        rom_memory[30830] = 3'b110;
        rom_memory[30831] = 3'b110;
        rom_memory[30832] = 3'b110;
        rom_memory[30833] = 3'b110;
        rom_memory[30834] = 3'b110;
        rom_memory[30835] = 3'b110;
        rom_memory[30836] = 3'b110;
        rom_memory[30837] = 3'b110;
        rom_memory[30838] = 3'b110;
        rom_memory[30839] = 3'b110;
        rom_memory[30840] = 3'b110;
        rom_memory[30841] = 3'b110;
        rom_memory[30842] = 3'b110;
        rom_memory[30843] = 3'b110;
        rom_memory[30844] = 3'b110;
        rom_memory[30845] = 3'b110;
        rom_memory[30846] = 3'b100;
        rom_memory[30847] = 3'b100;
        rom_memory[30848] = 3'b100;
        rom_memory[30849] = 3'b000;
        rom_memory[30850] = 3'b000;
        rom_memory[30851] = 3'b000;
        rom_memory[30852] = 3'b000;
        rom_memory[30853] = 3'b100;
        rom_memory[30854] = 3'b110;
        rom_memory[30855] = 3'b110;
        rom_memory[30856] = 3'b110;
        rom_memory[30857] = 3'b110;
        rom_memory[30858] = 3'b100;
        rom_memory[30859] = 3'b110;
        rom_memory[30860] = 3'b110;
        rom_memory[30861] = 3'b110;
        rom_memory[30862] = 3'b111;
        rom_memory[30863] = 3'b110;
        rom_memory[30864] = 3'b110;
        rom_memory[30865] = 3'b110;
        rom_memory[30866] = 3'b110;
        rom_memory[30867] = 3'b110;
        rom_memory[30868] = 3'b110;
        rom_memory[30869] = 3'b110;
        rom_memory[30870] = 3'b110;
        rom_memory[30871] = 3'b110;
        rom_memory[30872] = 3'b110;
        rom_memory[30873] = 3'b110;
        rom_memory[30874] = 3'b110;
        rom_memory[30875] = 3'b110;
        rom_memory[30876] = 3'b110;
        rom_memory[30877] = 3'b110;
        rom_memory[30878] = 3'b110;
        rom_memory[30879] = 3'b110;
        rom_memory[30880] = 3'b110;
        rom_memory[30881] = 3'b110;
        rom_memory[30882] = 3'b110;
        rom_memory[30883] = 3'b110;
        rom_memory[30884] = 3'b110;
        rom_memory[30885] = 3'b110;
        rom_memory[30886] = 3'b110;
        rom_memory[30887] = 3'b110;
        rom_memory[30888] = 3'b110;
        rom_memory[30889] = 3'b110;
        rom_memory[30890] = 3'b110;
        rom_memory[30891] = 3'b110;
        rom_memory[30892] = 3'b110;
        rom_memory[30893] = 3'b110;
        rom_memory[30894] = 3'b110;
        rom_memory[30895] = 3'b110;
        rom_memory[30896] = 3'b110;
        rom_memory[30897] = 3'b110;
        rom_memory[30898] = 3'b110;
        rom_memory[30899] = 3'b110;
        rom_memory[30900] = 3'b110;
        rom_memory[30901] = 3'b110;
        rom_memory[30902] = 3'b110;
        rom_memory[30903] = 3'b110;
        rom_memory[30904] = 3'b111;
        rom_memory[30905] = 3'b111;
        rom_memory[30906] = 3'b111;
        rom_memory[30907] = 3'b111;
        rom_memory[30908] = 3'b111;
        rom_memory[30909] = 3'b111;
        rom_memory[30910] = 3'b111;
        rom_memory[30911] = 3'b111;
        rom_memory[30912] = 3'b111;
        rom_memory[30913] = 3'b111;
        rom_memory[30914] = 3'b111;
        rom_memory[30915] = 3'b111;
        rom_memory[30916] = 3'b111;
        rom_memory[30917] = 3'b111;
        rom_memory[30918] = 3'b111;
        rom_memory[30919] = 3'b111;
        rom_memory[30920] = 3'b111;
        rom_memory[30921] = 3'b111;
        rom_memory[30922] = 3'b111;
        rom_memory[30923] = 3'b111;
        rom_memory[30924] = 3'b111;
        rom_memory[30925] = 3'b111;
        rom_memory[30926] = 3'b111;
        rom_memory[30927] = 3'b111;
        rom_memory[30928] = 3'b111;
        rom_memory[30929] = 3'b111;
        rom_memory[30930] = 3'b111;
        rom_memory[30931] = 3'b111;
        rom_memory[30932] = 3'b111;
        rom_memory[30933] = 3'b111;
        rom_memory[30934] = 3'b111;
        rom_memory[30935] = 3'b111;
        rom_memory[30936] = 3'b111;
        rom_memory[30937] = 3'b111;
        rom_memory[30938] = 3'b111;
        rom_memory[30939] = 3'b111;
        rom_memory[30940] = 3'b111;
        rom_memory[30941] = 3'b111;
        rom_memory[30942] = 3'b111;
        rom_memory[30943] = 3'b111;
        rom_memory[30944] = 3'b111;
        rom_memory[30945] = 3'b111;
        rom_memory[30946] = 3'b111;
        rom_memory[30947] = 3'b111;
        rom_memory[30948] = 3'b111;
        rom_memory[30949] = 3'b111;
        rom_memory[30950] = 3'b111;
        rom_memory[30951] = 3'b111;
        rom_memory[30952] = 3'b111;
        rom_memory[30953] = 3'b111;
        rom_memory[30954] = 3'b111;
        rom_memory[30955] = 3'b111;
        rom_memory[30956] = 3'b111;
        rom_memory[30957] = 3'b111;
        rom_memory[30958] = 3'b111;
        rom_memory[30959] = 3'b111;
        rom_memory[30960] = 3'b110;
        rom_memory[30961] = 3'b110;
        rom_memory[30962] = 3'b110;
        rom_memory[30963] = 3'b110;
        rom_memory[30964] = 3'b110;
        rom_memory[30965] = 3'b110;
        rom_memory[30966] = 3'b110;
        rom_memory[30967] = 3'b110;
        rom_memory[30968] = 3'b110;
        rom_memory[30969] = 3'b110;
        rom_memory[30970] = 3'b110;
        rom_memory[30971] = 3'b110;
        rom_memory[30972] = 3'b111;
        rom_memory[30973] = 3'b111;
        rom_memory[30974] = 3'b111;
        rom_memory[30975] = 3'b111;
        rom_memory[30976] = 3'b111;
        rom_memory[30977] = 3'b111;
        rom_memory[30978] = 3'b111;
        rom_memory[30979] = 3'b111;
        rom_memory[30980] = 3'b111;
        rom_memory[30981] = 3'b111;
        rom_memory[30982] = 3'b111;
        rom_memory[30983] = 3'b111;
        rom_memory[30984] = 3'b110;
        rom_memory[30985] = 3'b111;
        rom_memory[30986] = 3'b111;
        rom_memory[30987] = 3'b111;
        rom_memory[30988] = 3'b111;
        rom_memory[30989] = 3'b111;
        rom_memory[30990] = 3'b111;
        rom_memory[30991] = 3'b111;
        rom_memory[30992] = 3'b111;
        rom_memory[30993] = 3'b111;
        rom_memory[30994] = 3'b111;
        rom_memory[30995] = 3'b111;
        rom_memory[30996] = 3'b111;
        rom_memory[30997] = 3'b110;
        rom_memory[30998] = 3'b111;
        rom_memory[30999] = 3'b111;
        rom_memory[31000] = 3'b111;
        rom_memory[31001] = 3'b111;
        rom_memory[31002] = 3'b110;
        rom_memory[31003] = 3'b110;
        rom_memory[31004] = 3'b110;
        rom_memory[31005] = 3'b111;
        rom_memory[31006] = 3'b111;
        rom_memory[31007] = 3'b111;
        rom_memory[31008] = 3'b111;
        rom_memory[31009] = 3'b111;
        rom_memory[31010] = 3'b111;
        rom_memory[31011] = 3'b111;
        rom_memory[31012] = 3'b111;
        rom_memory[31013] = 3'b111;
        rom_memory[31014] = 3'b111;
        rom_memory[31015] = 3'b111;
        rom_memory[31016] = 3'b111;
        rom_memory[31017] = 3'b111;
        rom_memory[31018] = 3'b111;
        rom_memory[31019] = 3'b111;
        rom_memory[31020] = 3'b111;
        rom_memory[31021] = 3'b111;
        rom_memory[31022] = 3'b111;
        rom_memory[31023] = 3'b111;
        rom_memory[31024] = 3'b111;
        rom_memory[31025] = 3'b110;
        rom_memory[31026] = 3'b110;
        rom_memory[31027] = 3'b110;
        rom_memory[31028] = 3'b000;
        rom_memory[31029] = 3'b000;
        rom_memory[31030] = 3'b000;
        rom_memory[31031] = 3'b000;
        rom_memory[31032] = 3'b000;
        rom_memory[31033] = 3'b000;
        rom_memory[31034] = 3'b000;
        rom_memory[31035] = 3'b000;
        rom_memory[31036] = 3'b000;
        rom_memory[31037] = 3'b111;
        rom_memory[31038] = 3'b111;
        rom_memory[31039] = 3'b110;
        rom_memory[31040] = 3'b110;
        rom_memory[31041] = 3'b111;
        rom_memory[31042] = 3'b111;
        rom_memory[31043] = 3'b111;
        rom_memory[31044] = 3'b000;
        rom_memory[31045] = 3'b110;
        rom_memory[31046] = 3'b000;
        rom_memory[31047] = 3'b000;
        rom_memory[31048] = 3'b100;
        rom_memory[31049] = 3'b110;
        rom_memory[31050] = 3'b110;
        rom_memory[31051] = 3'b100;
        rom_memory[31052] = 3'b000;
        rom_memory[31053] = 3'b000;
        rom_memory[31054] = 3'b110;
        rom_memory[31055] = 3'b111;
        rom_memory[31056] = 3'b110;
        rom_memory[31057] = 3'b100;
        rom_memory[31058] = 3'b101;
        rom_memory[31059] = 3'b000;
        rom_memory[31060] = 3'b110;
        rom_memory[31061] = 3'b110;
        rom_memory[31062] = 3'b110;
        rom_memory[31063] = 3'b110;
        rom_memory[31064] = 3'b110;
        rom_memory[31065] = 3'b110;
        rom_memory[31066] = 3'b110;
        rom_memory[31067] = 3'b110;
        rom_memory[31068] = 3'b111;
        rom_memory[31069] = 3'b110;
        rom_memory[31070] = 3'b110;
        rom_memory[31071] = 3'b110;
        rom_memory[31072] = 3'b110;
        rom_memory[31073] = 3'b110;
        rom_memory[31074] = 3'b110;
        rom_memory[31075] = 3'b110;
        rom_memory[31076] = 3'b110;
        rom_memory[31077] = 3'b110;
        rom_memory[31078] = 3'b110;
        rom_memory[31079] = 3'b110;
        rom_memory[31080] = 3'b110;
        rom_memory[31081] = 3'b110;
        rom_memory[31082] = 3'b110;
        rom_memory[31083] = 3'b110;
        rom_memory[31084] = 3'b110;
        rom_memory[31085] = 3'b110;
        rom_memory[31086] = 3'b110;
        rom_memory[31087] = 3'b000;
        rom_memory[31088] = 3'b000;
        rom_memory[31089] = 3'b000;
        rom_memory[31090] = 3'b000;
        rom_memory[31091] = 3'b000;
        rom_memory[31092] = 3'b000;
        rom_memory[31093] = 3'b000;
        rom_memory[31094] = 3'b100;
        rom_memory[31095] = 3'b110;
        rom_memory[31096] = 3'b110;
        rom_memory[31097] = 3'b110;
        rom_memory[31098] = 3'b110;
        rom_memory[31099] = 3'b110;
        rom_memory[31100] = 3'b100;
        rom_memory[31101] = 3'b100;
        rom_memory[31102] = 3'b110;
        rom_memory[31103] = 3'b111;
        rom_memory[31104] = 3'b110;
        rom_memory[31105] = 3'b110;
        rom_memory[31106] = 3'b110;
        rom_memory[31107] = 3'b110;
        rom_memory[31108] = 3'b110;
        rom_memory[31109] = 3'b110;
        rom_memory[31110] = 3'b110;
        rom_memory[31111] = 3'b110;
        rom_memory[31112] = 3'b110;
        rom_memory[31113] = 3'b110;
        rom_memory[31114] = 3'b110;
        rom_memory[31115] = 3'b110;
        rom_memory[31116] = 3'b110;
        rom_memory[31117] = 3'b110;
        rom_memory[31118] = 3'b110;
        rom_memory[31119] = 3'b110;
        rom_memory[31120] = 3'b110;
        rom_memory[31121] = 3'b110;
        rom_memory[31122] = 3'b110;
        rom_memory[31123] = 3'b110;
        rom_memory[31124] = 3'b110;
        rom_memory[31125] = 3'b110;
        rom_memory[31126] = 3'b110;
        rom_memory[31127] = 3'b110;
        rom_memory[31128] = 3'b110;
        rom_memory[31129] = 3'b110;
        rom_memory[31130] = 3'b110;
        rom_memory[31131] = 3'b110;
        rom_memory[31132] = 3'b110;
        rom_memory[31133] = 3'b110;
        rom_memory[31134] = 3'b110;
        rom_memory[31135] = 3'b110;
        rom_memory[31136] = 3'b110;
        rom_memory[31137] = 3'b110;
        rom_memory[31138] = 3'b110;
        rom_memory[31139] = 3'b110;
        rom_memory[31140] = 3'b110;
        rom_memory[31141] = 3'b110;
        rom_memory[31142] = 3'b110;
        rom_memory[31143] = 3'b111;
        rom_memory[31144] = 3'b111;
        rom_memory[31145] = 3'b111;
        rom_memory[31146] = 3'b111;
        rom_memory[31147] = 3'b111;
        rom_memory[31148] = 3'b111;
        rom_memory[31149] = 3'b111;
        rom_memory[31150] = 3'b111;
        rom_memory[31151] = 3'b111;
        rom_memory[31152] = 3'b111;
        rom_memory[31153] = 3'b111;
        rom_memory[31154] = 3'b111;
        rom_memory[31155] = 3'b111;
        rom_memory[31156] = 3'b111;
        rom_memory[31157] = 3'b111;
        rom_memory[31158] = 3'b111;
        rom_memory[31159] = 3'b111;
        rom_memory[31160] = 3'b111;
        rom_memory[31161] = 3'b111;
        rom_memory[31162] = 3'b111;
        rom_memory[31163] = 3'b111;
        rom_memory[31164] = 3'b111;
        rom_memory[31165] = 3'b111;
        rom_memory[31166] = 3'b111;
        rom_memory[31167] = 3'b111;
        rom_memory[31168] = 3'b111;
        rom_memory[31169] = 3'b111;
        rom_memory[31170] = 3'b111;
        rom_memory[31171] = 3'b111;
        rom_memory[31172] = 3'b111;
        rom_memory[31173] = 3'b111;
        rom_memory[31174] = 3'b111;
        rom_memory[31175] = 3'b111;
        rom_memory[31176] = 3'b111;
        rom_memory[31177] = 3'b111;
        rom_memory[31178] = 3'b111;
        rom_memory[31179] = 3'b111;
        rom_memory[31180] = 3'b111;
        rom_memory[31181] = 3'b111;
        rom_memory[31182] = 3'b111;
        rom_memory[31183] = 3'b111;
        rom_memory[31184] = 3'b111;
        rom_memory[31185] = 3'b111;
        rom_memory[31186] = 3'b111;
        rom_memory[31187] = 3'b111;
        rom_memory[31188] = 3'b111;
        rom_memory[31189] = 3'b111;
        rom_memory[31190] = 3'b111;
        rom_memory[31191] = 3'b111;
        rom_memory[31192] = 3'b111;
        rom_memory[31193] = 3'b111;
        rom_memory[31194] = 3'b111;
        rom_memory[31195] = 3'b111;
        rom_memory[31196] = 3'b111;
        rom_memory[31197] = 3'b111;
        rom_memory[31198] = 3'b111;
        rom_memory[31199] = 3'b111;
        rom_memory[31200] = 3'b110;
        rom_memory[31201] = 3'b110;
        rom_memory[31202] = 3'b110;
        rom_memory[31203] = 3'b110;
        rom_memory[31204] = 3'b110;
        rom_memory[31205] = 3'b110;
        rom_memory[31206] = 3'b110;
        rom_memory[31207] = 3'b110;
        rom_memory[31208] = 3'b110;
        rom_memory[31209] = 3'b110;
        rom_memory[31210] = 3'b110;
        rom_memory[31211] = 3'b110;
        rom_memory[31212] = 3'b110;
        rom_memory[31213] = 3'b111;
        rom_memory[31214] = 3'b111;
        rom_memory[31215] = 3'b111;
        rom_memory[31216] = 3'b111;
        rom_memory[31217] = 3'b111;
        rom_memory[31218] = 3'b111;
        rom_memory[31219] = 3'b111;
        rom_memory[31220] = 3'b111;
        rom_memory[31221] = 3'b110;
        rom_memory[31222] = 3'b110;
        rom_memory[31223] = 3'b111;
        rom_memory[31224] = 3'b110;
        rom_memory[31225] = 3'b111;
        rom_memory[31226] = 3'b111;
        rom_memory[31227] = 3'b111;
        rom_memory[31228] = 3'b111;
        rom_memory[31229] = 3'b111;
        rom_memory[31230] = 3'b111;
        rom_memory[31231] = 3'b111;
        rom_memory[31232] = 3'b111;
        rom_memory[31233] = 3'b111;
        rom_memory[31234] = 3'b111;
        rom_memory[31235] = 3'b110;
        rom_memory[31236] = 3'b111;
        rom_memory[31237] = 3'b111;
        rom_memory[31238] = 3'b111;
        rom_memory[31239] = 3'b111;
        rom_memory[31240] = 3'b111;
        rom_memory[31241] = 3'b111;
        rom_memory[31242] = 3'b110;
        rom_memory[31243] = 3'b110;
        rom_memory[31244] = 3'b111;
        rom_memory[31245] = 3'b110;
        rom_memory[31246] = 3'b111;
        rom_memory[31247] = 3'b111;
        rom_memory[31248] = 3'b111;
        rom_memory[31249] = 3'b111;
        rom_memory[31250] = 3'b111;
        rom_memory[31251] = 3'b111;
        rom_memory[31252] = 3'b111;
        rom_memory[31253] = 3'b111;
        rom_memory[31254] = 3'b111;
        rom_memory[31255] = 3'b111;
        rom_memory[31256] = 3'b111;
        rom_memory[31257] = 3'b111;
        rom_memory[31258] = 3'b111;
        rom_memory[31259] = 3'b111;
        rom_memory[31260] = 3'b111;
        rom_memory[31261] = 3'b111;
        rom_memory[31262] = 3'b111;
        rom_memory[31263] = 3'b111;
        rom_memory[31264] = 3'b111;
        rom_memory[31265] = 3'b110;
        rom_memory[31266] = 3'b000;
        rom_memory[31267] = 3'b000;
        rom_memory[31268] = 3'b000;
        rom_memory[31269] = 3'b000;
        rom_memory[31270] = 3'b000;
        rom_memory[31271] = 3'b000;
        rom_memory[31272] = 3'b000;
        rom_memory[31273] = 3'b000;
        rom_memory[31274] = 3'b000;
        rom_memory[31275] = 3'b000;
        rom_memory[31276] = 3'b000;
        rom_memory[31277] = 3'b100;
        rom_memory[31278] = 3'b110;
        rom_memory[31279] = 3'b110;
        rom_memory[31280] = 3'b110;
        rom_memory[31281] = 3'b111;
        rom_memory[31282] = 3'b111;
        rom_memory[31283] = 3'b111;
        rom_memory[31284] = 3'b000;
        rom_memory[31285] = 3'b000;
        rom_memory[31286] = 3'b000;
        rom_memory[31287] = 3'b000;
        rom_memory[31288] = 3'b110;
        rom_memory[31289] = 3'b111;
        rom_memory[31290] = 3'b100;
        rom_memory[31291] = 3'b100;
        rom_memory[31292] = 3'b000;
        rom_memory[31293] = 3'b000;
        rom_memory[31294] = 3'b100;
        rom_memory[31295] = 3'b111;
        rom_memory[31296] = 3'b111;
        rom_memory[31297] = 3'b111;
        rom_memory[31298] = 3'b111;
        rom_memory[31299] = 3'b110;
        rom_memory[31300] = 3'b110;
        rom_memory[31301] = 3'b110;
        rom_memory[31302] = 3'b110;
        rom_memory[31303] = 3'b110;
        rom_memory[31304] = 3'b110;
        rom_memory[31305] = 3'b110;
        rom_memory[31306] = 3'b110;
        rom_memory[31307] = 3'b110;
        rom_memory[31308] = 3'b110;
        rom_memory[31309] = 3'b110;
        rom_memory[31310] = 3'b110;
        rom_memory[31311] = 3'b110;
        rom_memory[31312] = 3'b110;
        rom_memory[31313] = 3'b110;
        rom_memory[31314] = 3'b110;
        rom_memory[31315] = 3'b110;
        rom_memory[31316] = 3'b110;
        rom_memory[31317] = 3'b110;
        rom_memory[31318] = 3'b110;
        rom_memory[31319] = 3'b110;
        rom_memory[31320] = 3'b110;
        rom_memory[31321] = 3'b110;
        rom_memory[31322] = 3'b110;
        rom_memory[31323] = 3'b110;
        rom_memory[31324] = 3'b110;
        rom_memory[31325] = 3'b110;
        rom_memory[31326] = 3'b110;
        rom_memory[31327] = 3'b110;
        rom_memory[31328] = 3'b000;
        rom_memory[31329] = 3'b000;
        rom_memory[31330] = 3'b000;
        rom_memory[31331] = 3'b000;
        rom_memory[31332] = 3'b000;
        rom_memory[31333] = 3'b000;
        rom_memory[31334] = 3'b000;
        rom_memory[31335] = 3'b100;
        rom_memory[31336] = 3'b100;
        rom_memory[31337] = 3'b110;
        rom_memory[31338] = 3'b110;
        rom_memory[31339] = 3'b110;
        rom_memory[31340] = 3'b110;
        rom_memory[31341] = 3'b100;
        rom_memory[31342] = 3'b100;
        rom_memory[31343] = 3'b110;
        rom_memory[31344] = 3'b111;
        rom_memory[31345] = 3'b110;
        rom_memory[31346] = 3'b110;
        rom_memory[31347] = 3'b110;
        rom_memory[31348] = 3'b110;
        rom_memory[31349] = 3'b110;
        rom_memory[31350] = 3'b110;
        rom_memory[31351] = 3'b110;
        rom_memory[31352] = 3'b110;
        rom_memory[31353] = 3'b110;
        rom_memory[31354] = 3'b110;
        rom_memory[31355] = 3'b110;
        rom_memory[31356] = 3'b110;
        rom_memory[31357] = 3'b110;
        rom_memory[31358] = 3'b110;
        rom_memory[31359] = 3'b110;
        rom_memory[31360] = 3'b110;
        rom_memory[31361] = 3'b110;
        rom_memory[31362] = 3'b110;
        rom_memory[31363] = 3'b110;
        rom_memory[31364] = 3'b110;
        rom_memory[31365] = 3'b110;
        rom_memory[31366] = 3'b110;
        rom_memory[31367] = 3'b110;
        rom_memory[31368] = 3'b110;
        rom_memory[31369] = 3'b110;
        rom_memory[31370] = 3'b110;
        rom_memory[31371] = 3'b110;
        rom_memory[31372] = 3'b110;
        rom_memory[31373] = 3'b110;
        rom_memory[31374] = 3'b110;
        rom_memory[31375] = 3'b110;
        rom_memory[31376] = 3'b110;
        rom_memory[31377] = 3'b110;
        rom_memory[31378] = 3'b110;
        rom_memory[31379] = 3'b110;
        rom_memory[31380] = 3'b110;
        rom_memory[31381] = 3'b110;
        rom_memory[31382] = 3'b110;
        rom_memory[31383] = 3'b110;
        rom_memory[31384] = 3'b111;
        rom_memory[31385] = 3'b111;
        rom_memory[31386] = 3'b111;
        rom_memory[31387] = 3'b111;
        rom_memory[31388] = 3'b111;
        rom_memory[31389] = 3'b111;
        rom_memory[31390] = 3'b111;
        rom_memory[31391] = 3'b111;
        rom_memory[31392] = 3'b111;
        rom_memory[31393] = 3'b111;
        rom_memory[31394] = 3'b111;
        rom_memory[31395] = 3'b111;
        rom_memory[31396] = 3'b111;
        rom_memory[31397] = 3'b111;
        rom_memory[31398] = 3'b111;
        rom_memory[31399] = 3'b111;
        rom_memory[31400] = 3'b111;
        rom_memory[31401] = 3'b111;
        rom_memory[31402] = 3'b111;
        rom_memory[31403] = 3'b111;
        rom_memory[31404] = 3'b111;
        rom_memory[31405] = 3'b111;
        rom_memory[31406] = 3'b111;
        rom_memory[31407] = 3'b111;
        rom_memory[31408] = 3'b111;
        rom_memory[31409] = 3'b111;
        rom_memory[31410] = 3'b111;
        rom_memory[31411] = 3'b111;
        rom_memory[31412] = 3'b111;
        rom_memory[31413] = 3'b111;
        rom_memory[31414] = 3'b111;
        rom_memory[31415] = 3'b111;
        rom_memory[31416] = 3'b111;
        rom_memory[31417] = 3'b111;
        rom_memory[31418] = 3'b111;
        rom_memory[31419] = 3'b111;
        rom_memory[31420] = 3'b111;
        rom_memory[31421] = 3'b111;
        rom_memory[31422] = 3'b111;
        rom_memory[31423] = 3'b111;
        rom_memory[31424] = 3'b111;
        rom_memory[31425] = 3'b111;
        rom_memory[31426] = 3'b111;
        rom_memory[31427] = 3'b111;
        rom_memory[31428] = 3'b111;
        rom_memory[31429] = 3'b111;
        rom_memory[31430] = 3'b111;
        rom_memory[31431] = 3'b111;
        rom_memory[31432] = 3'b111;
        rom_memory[31433] = 3'b111;
        rom_memory[31434] = 3'b111;
        rom_memory[31435] = 3'b111;
        rom_memory[31436] = 3'b111;
        rom_memory[31437] = 3'b111;
        rom_memory[31438] = 3'b111;
        rom_memory[31439] = 3'b111;
        rom_memory[31440] = 3'b110;
        rom_memory[31441] = 3'b110;
        rom_memory[31442] = 3'b110;
        rom_memory[31443] = 3'b110;
        rom_memory[31444] = 3'b110;
        rom_memory[31445] = 3'b110;
        rom_memory[31446] = 3'b110;
        rom_memory[31447] = 3'b110;
        rom_memory[31448] = 3'b110;
        rom_memory[31449] = 3'b110;
        rom_memory[31450] = 3'b110;
        rom_memory[31451] = 3'b110;
        rom_memory[31452] = 3'b111;
        rom_memory[31453] = 3'b111;
        rom_memory[31454] = 3'b111;
        rom_memory[31455] = 3'b111;
        rom_memory[31456] = 3'b111;
        rom_memory[31457] = 3'b111;
        rom_memory[31458] = 3'b111;
        rom_memory[31459] = 3'b111;
        rom_memory[31460] = 3'b110;
        rom_memory[31461] = 3'b110;
        rom_memory[31462] = 3'b110;
        rom_memory[31463] = 3'b110;
        rom_memory[31464] = 3'b110;
        rom_memory[31465] = 3'b111;
        rom_memory[31466] = 3'b111;
        rom_memory[31467] = 3'b111;
        rom_memory[31468] = 3'b111;
        rom_memory[31469] = 3'b111;
        rom_memory[31470] = 3'b111;
        rom_memory[31471] = 3'b111;
        rom_memory[31472] = 3'b111;
        rom_memory[31473] = 3'b111;
        rom_memory[31474] = 3'b111;
        rom_memory[31475] = 3'b110;
        rom_memory[31476] = 3'b111;
        rom_memory[31477] = 3'b111;
        rom_memory[31478] = 3'b111;
        rom_memory[31479] = 3'b111;
        rom_memory[31480] = 3'b111;
        rom_memory[31481] = 3'b111;
        rom_memory[31482] = 3'b111;
        rom_memory[31483] = 3'b110;
        rom_memory[31484] = 3'b110;
        rom_memory[31485] = 3'b110;
        rom_memory[31486] = 3'b111;
        rom_memory[31487] = 3'b111;
        rom_memory[31488] = 3'b111;
        rom_memory[31489] = 3'b111;
        rom_memory[31490] = 3'b111;
        rom_memory[31491] = 3'b111;
        rom_memory[31492] = 3'b111;
        rom_memory[31493] = 3'b111;
        rom_memory[31494] = 3'b111;
        rom_memory[31495] = 3'b111;
        rom_memory[31496] = 3'b111;
        rom_memory[31497] = 3'b111;
        rom_memory[31498] = 3'b111;
        rom_memory[31499] = 3'b111;
        rom_memory[31500] = 3'b111;
        rom_memory[31501] = 3'b111;
        rom_memory[31502] = 3'b111;
        rom_memory[31503] = 3'b111;
        rom_memory[31504] = 3'b000;
        rom_memory[31505] = 3'b000;
        rom_memory[31506] = 3'b000;
        rom_memory[31507] = 3'b000;
        rom_memory[31508] = 3'b000;
        rom_memory[31509] = 3'b000;
        rom_memory[31510] = 3'b000;
        rom_memory[31511] = 3'b000;
        rom_memory[31512] = 3'b000;
        rom_memory[31513] = 3'b000;
        rom_memory[31514] = 3'b000;
        rom_memory[31515] = 3'b000;
        rom_memory[31516] = 3'b000;
        rom_memory[31517] = 3'b000;
        rom_memory[31518] = 3'b110;
        rom_memory[31519] = 3'b110;
        rom_memory[31520] = 3'b110;
        rom_memory[31521] = 3'b111;
        rom_memory[31522] = 3'b111;
        rom_memory[31523] = 3'b110;
        rom_memory[31524] = 3'b000;
        rom_memory[31525] = 3'b000;
        rom_memory[31526] = 3'b000;
        rom_memory[31527] = 3'b100;
        rom_memory[31528] = 3'b000;
        rom_memory[31529] = 3'b100;
        rom_memory[31530] = 3'b100;
        rom_memory[31531] = 3'b110;
        rom_memory[31532] = 3'b000;
        rom_memory[31533] = 3'b000;
        rom_memory[31534] = 3'b100;
        rom_memory[31535] = 3'b110;
        rom_memory[31536] = 3'b111;
        rom_memory[31537] = 3'b111;
        rom_memory[31538] = 3'b111;
        rom_memory[31539] = 3'b111;
        rom_memory[31540] = 3'b110;
        rom_memory[31541] = 3'b110;
        rom_memory[31542] = 3'b110;
        rom_memory[31543] = 3'b110;
        rom_memory[31544] = 3'b110;
        rom_memory[31545] = 3'b110;
        rom_memory[31546] = 3'b110;
        rom_memory[31547] = 3'b110;
        rom_memory[31548] = 3'b110;
        rom_memory[31549] = 3'b110;
        rom_memory[31550] = 3'b110;
        rom_memory[31551] = 3'b110;
        rom_memory[31552] = 3'b110;
        rom_memory[31553] = 3'b110;
        rom_memory[31554] = 3'b110;
        rom_memory[31555] = 3'b110;
        rom_memory[31556] = 3'b110;
        rom_memory[31557] = 3'b110;
        rom_memory[31558] = 3'b110;
        rom_memory[31559] = 3'b110;
        rom_memory[31560] = 3'b110;
        rom_memory[31561] = 3'b110;
        rom_memory[31562] = 3'b110;
        rom_memory[31563] = 3'b110;
        rom_memory[31564] = 3'b110;
        rom_memory[31565] = 3'b110;
        rom_memory[31566] = 3'b110;
        rom_memory[31567] = 3'b110;
        rom_memory[31568] = 3'b110;
        rom_memory[31569] = 3'b000;
        rom_memory[31570] = 3'b000;
        rom_memory[31571] = 3'b000;
        rom_memory[31572] = 3'b000;
        rom_memory[31573] = 3'b000;
        rom_memory[31574] = 3'b000;
        rom_memory[31575] = 3'b000;
        rom_memory[31576] = 3'b000;
        rom_memory[31577] = 3'b100;
        rom_memory[31578] = 3'b110;
        rom_memory[31579] = 3'b110;
        rom_memory[31580] = 3'b110;
        rom_memory[31581] = 3'b100;
        rom_memory[31582] = 3'b100;
        rom_memory[31583] = 3'b100;
        rom_memory[31584] = 3'b110;
        rom_memory[31585] = 3'b111;
        rom_memory[31586] = 3'b110;
        rom_memory[31587] = 3'b110;
        rom_memory[31588] = 3'b110;
        rom_memory[31589] = 3'b110;
        rom_memory[31590] = 3'b110;
        rom_memory[31591] = 3'b110;
        rom_memory[31592] = 3'b110;
        rom_memory[31593] = 3'b110;
        rom_memory[31594] = 3'b110;
        rom_memory[31595] = 3'b110;
        rom_memory[31596] = 3'b110;
        rom_memory[31597] = 3'b110;
        rom_memory[31598] = 3'b110;
        rom_memory[31599] = 3'b110;
        rom_memory[31600] = 3'b110;
        rom_memory[31601] = 3'b110;
        rom_memory[31602] = 3'b110;
        rom_memory[31603] = 3'b110;
        rom_memory[31604] = 3'b110;
        rom_memory[31605] = 3'b110;
        rom_memory[31606] = 3'b110;
        rom_memory[31607] = 3'b110;
        rom_memory[31608] = 3'b110;
        rom_memory[31609] = 3'b110;
        rom_memory[31610] = 3'b110;
        rom_memory[31611] = 3'b110;
        rom_memory[31612] = 3'b110;
        rom_memory[31613] = 3'b110;
        rom_memory[31614] = 3'b110;
        rom_memory[31615] = 3'b110;
        rom_memory[31616] = 3'b110;
        rom_memory[31617] = 3'b110;
        rom_memory[31618] = 3'b110;
        rom_memory[31619] = 3'b110;
        rom_memory[31620] = 3'b110;
        rom_memory[31621] = 3'b111;
        rom_memory[31622] = 3'b110;
        rom_memory[31623] = 3'b111;
        rom_memory[31624] = 3'b111;
        rom_memory[31625] = 3'b111;
        rom_memory[31626] = 3'b111;
        rom_memory[31627] = 3'b111;
        rom_memory[31628] = 3'b111;
        rom_memory[31629] = 3'b111;
        rom_memory[31630] = 3'b111;
        rom_memory[31631] = 3'b111;
        rom_memory[31632] = 3'b111;
        rom_memory[31633] = 3'b111;
        rom_memory[31634] = 3'b111;
        rom_memory[31635] = 3'b111;
        rom_memory[31636] = 3'b111;
        rom_memory[31637] = 3'b111;
        rom_memory[31638] = 3'b111;
        rom_memory[31639] = 3'b111;
        rom_memory[31640] = 3'b111;
        rom_memory[31641] = 3'b111;
        rom_memory[31642] = 3'b111;
        rom_memory[31643] = 3'b111;
        rom_memory[31644] = 3'b111;
        rom_memory[31645] = 3'b111;
        rom_memory[31646] = 3'b111;
        rom_memory[31647] = 3'b111;
        rom_memory[31648] = 3'b111;
        rom_memory[31649] = 3'b111;
        rom_memory[31650] = 3'b111;
        rom_memory[31651] = 3'b111;
        rom_memory[31652] = 3'b111;
        rom_memory[31653] = 3'b111;
        rom_memory[31654] = 3'b111;
        rom_memory[31655] = 3'b111;
        rom_memory[31656] = 3'b111;
        rom_memory[31657] = 3'b111;
        rom_memory[31658] = 3'b111;
        rom_memory[31659] = 3'b111;
        rom_memory[31660] = 3'b111;
        rom_memory[31661] = 3'b111;
        rom_memory[31662] = 3'b111;
        rom_memory[31663] = 3'b111;
        rom_memory[31664] = 3'b111;
        rom_memory[31665] = 3'b111;
        rom_memory[31666] = 3'b111;
        rom_memory[31667] = 3'b111;
        rom_memory[31668] = 3'b111;
        rom_memory[31669] = 3'b111;
        rom_memory[31670] = 3'b111;
        rom_memory[31671] = 3'b111;
        rom_memory[31672] = 3'b111;
        rom_memory[31673] = 3'b111;
        rom_memory[31674] = 3'b111;
        rom_memory[31675] = 3'b111;
        rom_memory[31676] = 3'b111;
        rom_memory[31677] = 3'b111;
        rom_memory[31678] = 3'b111;
        rom_memory[31679] = 3'b111;
        rom_memory[31680] = 3'b110;
        rom_memory[31681] = 3'b110;
        rom_memory[31682] = 3'b110;
        rom_memory[31683] = 3'b110;
        rom_memory[31684] = 3'b110;
        rom_memory[31685] = 3'b110;
        rom_memory[31686] = 3'b110;
        rom_memory[31687] = 3'b110;
        rom_memory[31688] = 3'b110;
        rom_memory[31689] = 3'b110;
        rom_memory[31690] = 3'b111;
        rom_memory[31691] = 3'b111;
        rom_memory[31692] = 3'b111;
        rom_memory[31693] = 3'b111;
        rom_memory[31694] = 3'b111;
        rom_memory[31695] = 3'b111;
        rom_memory[31696] = 3'b111;
        rom_memory[31697] = 3'b111;
        rom_memory[31698] = 3'b111;
        rom_memory[31699] = 3'b111;
        rom_memory[31700] = 3'b110;
        rom_memory[31701] = 3'b110;
        rom_memory[31702] = 3'b110;
        rom_memory[31703] = 3'b110;
        rom_memory[31704] = 3'b110;
        rom_memory[31705] = 3'b110;
        rom_memory[31706] = 3'b111;
        rom_memory[31707] = 3'b111;
        rom_memory[31708] = 3'b111;
        rom_memory[31709] = 3'b111;
        rom_memory[31710] = 3'b111;
        rom_memory[31711] = 3'b111;
        rom_memory[31712] = 3'b111;
        rom_memory[31713] = 3'b111;
        rom_memory[31714] = 3'b111;
        rom_memory[31715] = 3'b110;
        rom_memory[31716] = 3'b110;
        rom_memory[31717] = 3'b111;
        rom_memory[31718] = 3'b111;
        rom_memory[31719] = 3'b111;
        rom_memory[31720] = 3'b111;
        rom_memory[31721] = 3'b111;
        rom_memory[31722] = 3'b111;
        rom_memory[31723] = 3'b110;
        rom_memory[31724] = 3'b110;
        rom_memory[31725] = 3'b110;
        rom_memory[31726] = 3'b111;
        rom_memory[31727] = 3'b111;
        rom_memory[31728] = 3'b111;
        rom_memory[31729] = 3'b111;
        rom_memory[31730] = 3'b111;
        rom_memory[31731] = 3'b111;
        rom_memory[31732] = 3'b111;
        rom_memory[31733] = 3'b111;
        rom_memory[31734] = 3'b111;
        rom_memory[31735] = 3'b111;
        rom_memory[31736] = 3'b111;
        rom_memory[31737] = 3'b111;
        rom_memory[31738] = 3'b111;
        rom_memory[31739] = 3'b111;
        rom_memory[31740] = 3'b111;
        rom_memory[31741] = 3'b111;
        rom_memory[31742] = 3'b111;
        rom_memory[31743] = 3'b001;
        rom_memory[31744] = 3'b000;
        rom_memory[31745] = 3'b000;
        rom_memory[31746] = 3'b000;
        rom_memory[31747] = 3'b000;
        rom_memory[31748] = 3'b000;
        rom_memory[31749] = 3'b000;
        rom_memory[31750] = 3'b000;
        rom_memory[31751] = 3'b000;
        rom_memory[31752] = 3'b000;
        rom_memory[31753] = 3'b000;
        rom_memory[31754] = 3'b000;
        rom_memory[31755] = 3'b000;
        rom_memory[31756] = 3'b110;
        rom_memory[31757] = 3'b000;
        rom_memory[31758] = 3'b110;
        rom_memory[31759] = 3'b110;
        rom_memory[31760] = 3'b110;
        rom_memory[31761] = 3'b110;
        rom_memory[31762] = 3'b111;
        rom_memory[31763] = 3'b111;
        rom_memory[31764] = 3'b110;
        rom_memory[31765] = 3'b000;
        rom_memory[31766] = 3'b000;
        rom_memory[31767] = 3'b000;
        rom_memory[31768] = 3'b000;
        rom_memory[31769] = 3'b000;
        rom_memory[31770] = 3'b110;
        rom_memory[31771] = 3'b110;
        rom_memory[31772] = 3'b100;
        rom_memory[31773] = 3'b110;
        rom_memory[31774] = 3'b111;
        rom_memory[31775] = 3'b111;
        rom_memory[31776] = 3'b000;
        rom_memory[31777] = 3'b000;
        rom_memory[31778] = 3'b111;
        rom_memory[31779] = 3'b111;
        rom_memory[31780] = 3'b110;
        rom_memory[31781] = 3'b110;
        rom_memory[31782] = 3'b110;
        rom_memory[31783] = 3'b110;
        rom_memory[31784] = 3'b110;
        rom_memory[31785] = 3'b110;
        rom_memory[31786] = 3'b110;
        rom_memory[31787] = 3'b110;
        rom_memory[31788] = 3'b110;
        rom_memory[31789] = 3'b110;
        rom_memory[31790] = 3'b110;
        rom_memory[31791] = 3'b110;
        rom_memory[31792] = 3'b110;
        rom_memory[31793] = 3'b110;
        rom_memory[31794] = 3'b110;
        rom_memory[31795] = 3'b110;
        rom_memory[31796] = 3'b110;
        rom_memory[31797] = 3'b110;
        rom_memory[31798] = 3'b110;
        rom_memory[31799] = 3'b110;
        rom_memory[31800] = 3'b110;
        rom_memory[31801] = 3'b110;
        rom_memory[31802] = 3'b110;
        rom_memory[31803] = 3'b110;
        rom_memory[31804] = 3'b110;
        rom_memory[31805] = 3'b110;
        rom_memory[31806] = 3'b110;
        rom_memory[31807] = 3'b110;
        rom_memory[31808] = 3'b110;
        rom_memory[31809] = 3'b110;
        rom_memory[31810] = 3'b000;
        rom_memory[31811] = 3'b000;
        rom_memory[31812] = 3'b000;
        rom_memory[31813] = 3'b000;
        rom_memory[31814] = 3'b000;
        rom_memory[31815] = 3'b000;
        rom_memory[31816] = 3'b000;
        rom_memory[31817] = 3'b000;
        rom_memory[31818] = 3'b000;
        rom_memory[31819] = 3'b100;
        rom_memory[31820] = 3'b110;
        rom_memory[31821] = 3'b110;
        rom_memory[31822] = 3'b100;
        rom_memory[31823] = 3'b000;
        rom_memory[31824] = 3'b100;
        rom_memory[31825] = 3'b110;
        rom_memory[31826] = 3'b111;
        rom_memory[31827] = 3'b110;
        rom_memory[31828] = 3'b110;
        rom_memory[31829] = 3'b110;
        rom_memory[31830] = 3'b110;
        rom_memory[31831] = 3'b110;
        rom_memory[31832] = 3'b110;
        rom_memory[31833] = 3'b110;
        rom_memory[31834] = 3'b110;
        rom_memory[31835] = 3'b110;
        rom_memory[31836] = 3'b110;
        rom_memory[31837] = 3'b110;
        rom_memory[31838] = 3'b110;
        rom_memory[31839] = 3'b110;
        rom_memory[31840] = 3'b110;
        rom_memory[31841] = 3'b110;
        rom_memory[31842] = 3'b110;
        rom_memory[31843] = 3'b110;
        rom_memory[31844] = 3'b110;
        rom_memory[31845] = 3'b110;
        rom_memory[31846] = 3'b110;
        rom_memory[31847] = 3'b110;
        rom_memory[31848] = 3'b110;
        rom_memory[31849] = 3'b110;
        rom_memory[31850] = 3'b110;
        rom_memory[31851] = 3'b110;
        rom_memory[31852] = 3'b110;
        rom_memory[31853] = 3'b110;
        rom_memory[31854] = 3'b110;
        rom_memory[31855] = 3'b110;
        rom_memory[31856] = 3'b110;
        rom_memory[31857] = 3'b110;
        rom_memory[31858] = 3'b110;
        rom_memory[31859] = 3'b110;
        rom_memory[31860] = 3'b110;
        rom_memory[31861] = 3'b110;
        rom_memory[31862] = 3'b110;
        rom_memory[31863] = 3'b111;
        rom_memory[31864] = 3'b111;
        rom_memory[31865] = 3'b111;
        rom_memory[31866] = 3'b111;
        rom_memory[31867] = 3'b111;
        rom_memory[31868] = 3'b111;
        rom_memory[31869] = 3'b111;
        rom_memory[31870] = 3'b111;
        rom_memory[31871] = 3'b111;
        rom_memory[31872] = 3'b111;
        rom_memory[31873] = 3'b111;
        rom_memory[31874] = 3'b111;
        rom_memory[31875] = 3'b111;
        rom_memory[31876] = 3'b111;
        rom_memory[31877] = 3'b111;
        rom_memory[31878] = 3'b111;
        rom_memory[31879] = 3'b111;
        rom_memory[31880] = 3'b111;
        rom_memory[31881] = 3'b111;
        rom_memory[31882] = 3'b111;
        rom_memory[31883] = 3'b111;
        rom_memory[31884] = 3'b111;
        rom_memory[31885] = 3'b111;
        rom_memory[31886] = 3'b111;
        rom_memory[31887] = 3'b111;
        rom_memory[31888] = 3'b111;
        rom_memory[31889] = 3'b111;
        rom_memory[31890] = 3'b111;
        rom_memory[31891] = 3'b111;
        rom_memory[31892] = 3'b111;
        rom_memory[31893] = 3'b111;
        rom_memory[31894] = 3'b111;
        rom_memory[31895] = 3'b111;
        rom_memory[31896] = 3'b111;
        rom_memory[31897] = 3'b111;
        rom_memory[31898] = 3'b111;
        rom_memory[31899] = 3'b111;
        rom_memory[31900] = 3'b111;
        rom_memory[31901] = 3'b111;
        rom_memory[31902] = 3'b111;
        rom_memory[31903] = 3'b111;
        rom_memory[31904] = 3'b111;
        rom_memory[31905] = 3'b111;
        rom_memory[31906] = 3'b111;
        rom_memory[31907] = 3'b111;
        rom_memory[31908] = 3'b111;
        rom_memory[31909] = 3'b111;
        rom_memory[31910] = 3'b111;
        rom_memory[31911] = 3'b111;
        rom_memory[31912] = 3'b111;
        rom_memory[31913] = 3'b111;
        rom_memory[31914] = 3'b111;
        rom_memory[31915] = 3'b111;
        rom_memory[31916] = 3'b111;
        rom_memory[31917] = 3'b111;
        rom_memory[31918] = 3'b111;
        rom_memory[31919] = 3'b111;
        rom_memory[31920] = 3'b110;
        rom_memory[31921] = 3'b110;
        rom_memory[31922] = 3'b110;
        rom_memory[31923] = 3'b110;
        rom_memory[31924] = 3'b110;
        rom_memory[31925] = 3'b110;
        rom_memory[31926] = 3'b110;
        rom_memory[31927] = 3'b110;
        rom_memory[31928] = 3'b110;
        rom_memory[31929] = 3'b111;
        rom_memory[31930] = 3'b111;
        rom_memory[31931] = 3'b111;
        rom_memory[31932] = 3'b111;
        rom_memory[31933] = 3'b111;
        rom_memory[31934] = 3'b111;
        rom_memory[31935] = 3'b111;
        rom_memory[31936] = 3'b111;
        rom_memory[31937] = 3'b111;
        rom_memory[31938] = 3'b111;
        rom_memory[31939] = 3'b111;
        rom_memory[31940] = 3'b110;
        rom_memory[31941] = 3'b110;
        rom_memory[31942] = 3'b110;
        rom_memory[31943] = 3'b110;
        rom_memory[31944] = 3'b110;
        rom_memory[31945] = 3'b110;
        rom_memory[31946] = 3'b111;
        rom_memory[31947] = 3'b111;
        rom_memory[31948] = 3'b111;
        rom_memory[31949] = 3'b111;
        rom_memory[31950] = 3'b111;
        rom_memory[31951] = 3'b111;
        rom_memory[31952] = 3'b111;
        rom_memory[31953] = 3'b111;
        rom_memory[31954] = 3'b111;
        rom_memory[31955] = 3'b110;
        rom_memory[31956] = 3'b110;
        rom_memory[31957] = 3'b111;
        rom_memory[31958] = 3'b111;
        rom_memory[31959] = 3'b111;
        rom_memory[31960] = 3'b111;
        rom_memory[31961] = 3'b111;
        rom_memory[31962] = 3'b110;
        rom_memory[31963] = 3'b110;
        rom_memory[31964] = 3'b110;
        rom_memory[31965] = 3'b110;
        rom_memory[31966] = 3'b111;
        rom_memory[31967] = 3'b111;
        rom_memory[31968] = 3'b111;
        rom_memory[31969] = 3'b111;
        rom_memory[31970] = 3'b111;
        rom_memory[31971] = 3'b111;
        rom_memory[31972] = 3'b111;
        rom_memory[31973] = 3'b111;
        rom_memory[31974] = 3'b111;
        rom_memory[31975] = 3'b111;
        rom_memory[31976] = 3'b111;
        rom_memory[31977] = 3'b111;
        rom_memory[31978] = 3'b111;
        rom_memory[31979] = 3'b111;
        rom_memory[31980] = 3'b111;
        rom_memory[31981] = 3'b111;
        rom_memory[31982] = 3'b111;
        rom_memory[31983] = 3'b000;
        rom_memory[31984] = 3'b000;
        rom_memory[31985] = 3'b000;
        rom_memory[31986] = 3'b000;
        rom_memory[31987] = 3'b000;
        rom_memory[31988] = 3'b000;
        rom_memory[31989] = 3'b000;
        rom_memory[31990] = 3'b000;
        rom_memory[31991] = 3'b000;
        rom_memory[31992] = 3'b000;
        rom_memory[31993] = 3'b000;
        rom_memory[31994] = 3'b000;
        rom_memory[31995] = 3'b110;
        rom_memory[31996] = 3'b111;
        rom_memory[31997] = 3'b111;
        rom_memory[31998] = 3'b100;
        rom_memory[31999] = 3'b110;
        rom_memory[32000] = 3'b110;
        rom_memory[32001] = 3'b110;
        rom_memory[32002] = 3'b111;
        rom_memory[32003] = 3'b110;
        rom_memory[32004] = 3'b111;
        rom_memory[32005] = 3'b111;
        rom_memory[32006] = 3'b000;
        rom_memory[32007] = 3'b000;
        rom_memory[32008] = 3'b000;
        rom_memory[32009] = 3'b100;
        rom_memory[32010] = 3'b100;
        rom_memory[32011] = 3'b100;
        rom_memory[32012] = 3'b000;
        rom_memory[32013] = 3'b100;
        rom_memory[32014] = 3'b111;
        rom_memory[32015] = 3'b111;
        rom_memory[32016] = 3'b111;
        rom_memory[32017] = 3'b000;
        rom_memory[32018] = 3'b111;
        rom_memory[32019] = 3'b111;
        rom_memory[32020] = 3'b111;
        rom_memory[32021] = 3'b110;
        rom_memory[32022] = 3'b110;
        rom_memory[32023] = 3'b110;
        rom_memory[32024] = 3'b110;
        rom_memory[32025] = 3'b110;
        rom_memory[32026] = 3'b110;
        rom_memory[32027] = 3'b110;
        rom_memory[32028] = 3'b110;
        rom_memory[32029] = 3'b110;
        rom_memory[32030] = 3'b110;
        rom_memory[32031] = 3'b110;
        rom_memory[32032] = 3'b110;
        rom_memory[32033] = 3'b110;
        rom_memory[32034] = 3'b110;
        rom_memory[32035] = 3'b110;
        rom_memory[32036] = 3'b110;
        rom_memory[32037] = 3'b110;
        rom_memory[32038] = 3'b110;
        rom_memory[32039] = 3'b110;
        rom_memory[32040] = 3'b110;
        rom_memory[32041] = 3'b110;
        rom_memory[32042] = 3'b110;
        rom_memory[32043] = 3'b110;
        rom_memory[32044] = 3'b110;
        rom_memory[32045] = 3'b110;
        rom_memory[32046] = 3'b110;
        rom_memory[32047] = 3'b110;
        rom_memory[32048] = 3'b110;
        rom_memory[32049] = 3'b110;
        rom_memory[32050] = 3'b111;
        rom_memory[32051] = 3'b100;
        rom_memory[32052] = 3'b000;
        rom_memory[32053] = 3'b000;
        rom_memory[32054] = 3'b000;
        rom_memory[32055] = 3'b000;
        rom_memory[32056] = 3'b000;
        rom_memory[32057] = 3'b000;
        rom_memory[32058] = 3'b000;
        rom_memory[32059] = 3'b000;
        rom_memory[32060] = 3'b100;
        rom_memory[32061] = 3'b110;
        rom_memory[32062] = 3'b110;
        rom_memory[32063] = 3'b100;
        rom_memory[32064] = 3'b000;
        rom_memory[32065] = 3'b100;
        rom_memory[32066] = 3'b110;
        rom_memory[32067] = 3'b111;
        rom_memory[32068] = 3'b110;
        rom_memory[32069] = 3'b110;
        rom_memory[32070] = 3'b110;
        rom_memory[32071] = 3'b110;
        rom_memory[32072] = 3'b110;
        rom_memory[32073] = 3'b110;
        rom_memory[32074] = 3'b110;
        rom_memory[32075] = 3'b110;
        rom_memory[32076] = 3'b110;
        rom_memory[32077] = 3'b110;
        rom_memory[32078] = 3'b110;
        rom_memory[32079] = 3'b110;
        rom_memory[32080] = 3'b110;
        rom_memory[32081] = 3'b110;
        rom_memory[32082] = 3'b110;
        rom_memory[32083] = 3'b110;
        rom_memory[32084] = 3'b110;
        rom_memory[32085] = 3'b110;
        rom_memory[32086] = 3'b110;
        rom_memory[32087] = 3'b110;
        rom_memory[32088] = 3'b110;
        rom_memory[32089] = 3'b110;
        rom_memory[32090] = 3'b110;
        rom_memory[32091] = 3'b110;
        rom_memory[32092] = 3'b110;
        rom_memory[32093] = 3'b110;
        rom_memory[32094] = 3'b110;
        rom_memory[32095] = 3'b110;
        rom_memory[32096] = 3'b110;
        rom_memory[32097] = 3'b110;
        rom_memory[32098] = 3'b110;
        rom_memory[32099] = 3'b110;
        rom_memory[32100] = 3'b110;
        rom_memory[32101] = 3'b110;
        rom_memory[32102] = 3'b110;
        rom_memory[32103] = 3'b111;
        rom_memory[32104] = 3'b111;
        rom_memory[32105] = 3'b111;
        rom_memory[32106] = 3'b111;
        rom_memory[32107] = 3'b111;
        rom_memory[32108] = 3'b111;
        rom_memory[32109] = 3'b111;
        rom_memory[32110] = 3'b111;
        rom_memory[32111] = 3'b111;
        rom_memory[32112] = 3'b111;
        rom_memory[32113] = 3'b111;
        rom_memory[32114] = 3'b111;
        rom_memory[32115] = 3'b111;
        rom_memory[32116] = 3'b111;
        rom_memory[32117] = 3'b111;
        rom_memory[32118] = 3'b111;
        rom_memory[32119] = 3'b111;
        rom_memory[32120] = 3'b111;
        rom_memory[32121] = 3'b111;
        rom_memory[32122] = 3'b111;
        rom_memory[32123] = 3'b111;
        rom_memory[32124] = 3'b111;
        rom_memory[32125] = 3'b111;
        rom_memory[32126] = 3'b111;
        rom_memory[32127] = 3'b111;
        rom_memory[32128] = 3'b111;
        rom_memory[32129] = 3'b111;
        rom_memory[32130] = 3'b111;
        rom_memory[32131] = 3'b111;
        rom_memory[32132] = 3'b111;
        rom_memory[32133] = 3'b111;
        rom_memory[32134] = 3'b111;
        rom_memory[32135] = 3'b111;
        rom_memory[32136] = 3'b111;
        rom_memory[32137] = 3'b111;
        rom_memory[32138] = 3'b111;
        rom_memory[32139] = 3'b111;
        rom_memory[32140] = 3'b111;
        rom_memory[32141] = 3'b111;
        rom_memory[32142] = 3'b111;
        rom_memory[32143] = 3'b111;
        rom_memory[32144] = 3'b111;
        rom_memory[32145] = 3'b111;
        rom_memory[32146] = 3'b111;
        rom_memory[32147] = 3'b111;
        rom_memory[32148] = 3'b111;
        rom_memory[32149] = 3'b111;
        rom_memory[32150] = 3'b111;
        rom_memory[32151] = 3'b111;
        rom_memory[32152] = 3'b111;
        rom_memory[32153] = 3'b111;
        rom_memory[32154] = 3'b111;
        rom_memory[32155] = 3'b111;
        rom_memory[32156] = 3'b111;
        rom_memory[32157] = 3'b111;
        rom_memory[32158] = 3'b111;
        rom_memory[32159] = 3'b111;
        rom_memory[32160] = 3'b110;
        rom_memory[32161] = 3'b110;
        rom_memory[32162] = 3'b110;
        rom_memory[32163] = 3'b110;
        rom_memory[32164] = 3'b110;
        rom_memory[32165] = 3'b110;
        rom_memory[32166] = 3'b110;
        rom_memory[32167] = 3'b110;
        rom_memory[32168] = 3'b110;
        rom_memory[32169] = 3'b111;
        rom_memory[32170] = 3'b111;
        rom_memory[32171] = 3'b111;
        rom_memory[32172] = 3'b111;
        rom_memory[32173] = 3'b111;
        rom_memory[32174] = 3'b111;
        rom_memory[32175] = 3'b111;
        rom_memory[32176] = 3'b111;
        rom_memory[32177] = 3'b111;
        rom_memory[32178] = 3'b111;
        rom_memory[32179] = 3'b111;
        rom_memory[32180] = 3'b110;
        rom_memory[32181] = 3'b110;
        rom_memory[32182] = 3'b110;
        rom_memory[32183] = 3'b110;
        rom_memory[32184] = 3'b110;
        rom_memory[32185] = 3'b110;
        rom_memory[32186] = 3'b111;
        rom_memory[32187] = 3'b111;
        rom_memory[32188] = 3'b111;
        rom_memory[32189] = 3'b111;
        rom_memory[32190] = 3'b111;
        rom_memory[32191] = 3'b111;
        rom_memory[32192] = 3'b111;
        rom_memory[32193] = 3'b111;
        rom_memory[32194] = 3'b111;
        rom_memory[32195] = 3'b111;
        rom_memory[32196] = 3'b110;
        rom_memory[32197] = 3'b111;
        rom_memory[32198] = 3'b111;
        rom_memory[32199] = 3'b111;
        rom_memory[32200] = 3'b111;
        rom_memory[32201] = 3'b110;
        rom_memory[32202] = 3'b110;
        rom_memory[32203] = 3'b110;
        rom_memory[32204] = 3'b110;
        rom_memory[32205] = 3'b110;
        rom_memory[32206] = 3'b111;
        rom_memory[32207] = 3'b111;
        rom_memory[32208] = 3'b111;
        rom_memory[32209] = 3'b111;
        rom_memory[32210] = 3'b111;
        rom_memory[32211] = 3'b111;
        rom_memory[32212] = 3'b111;
        rom_memory[32213] = 3'b111;
        rom_memory[32214] = 3'b111;
        rom_memory[32215] = 3'b111;
        rom_memory[32216] = 3'b111;
        rom_memory[32217] = 3'b111;
        rom_memory[32218] = 3'b111;
        rom_memory[32219] = 3'b111;
        rom_memory[32220] = 3'b111;
        rom_memory[32221] = 3'b111;
        rom_memory[32222] = 3'b000;
        rom_memory[32223] = 3'b000;
        rom_memory[32224] = 3'b000;
        rom_memory[32225] = 3'b000;
        rom_memory[32226] = 3'b000;
        rom_memory[32227] = 3'b000;
        rom_memory[32228] = 3'b000;
        rom_memory[32229] = 3'b000;
        rom_memory[32230] = 3'b000;
        rom_memory[32231] = 3'b000;
        rom_memory[32232] = 3'b000;
        rom_memory[32233] = 3'b000;
        rom_memory[32234] = 3'b111;
        rom_memory[32235] = 3'b111;
        rom_memory[32236] = 3'b111;
        rom_memory[32237] = 3'b111;
        rom_memory[32238] = 3'b110;
        rom_memory[32239] = 3'b110;
        rom_memory[32240] = 3'b110;
        rom_memory[32241] = 3'b110;
        rom_memory[32242] = 3'b110;
        rom_memory[32243] = 3'b110;
        rom_memory[32244] = 3'b110;
        rom_memory[32245] = 3'b111;
        rom_memory[32246] = 3'b111;
        rom_memory[32247] = 3'b000;
        rom_memory[32248] = 3'b111;
        rom_memory[32249] = 3'b111;
        rom_memory[32250] = 3'b100;
        rom_memory[32251] = 3'b000;
        rom_memory[32252] = 3'b000;
        rom_memory[32253] = 3'b111;
        rom_memory[32254] = 3'b111;
        rom_memory[32255] = 3'b100;
        rom_memory[32256] = 3'b100;
        rom_memory[32257] = 3'b111;
        rom_memory[32258] = 3'b111;
        rom_memory[32259] = 3'b111;
        rom_memory[32260] = 3'b110;
        rom_memory[32261] = 3'b110;
        rom_memory[32262] = 3'b110;
        rom_memory[32263] = 3'b110;
        rom_memory[32264] = 3'b110;
        rom_memory[32265] = 3'b110;
        rom_memory[32266] = 3'b110;
        rom_memory[32267] = 3'b110;
        rom_memory[32268] = 3'b110;
        rom_memory[32269] = 3'b110;
        rom_memory[32270] = 3'b110;
        rom_memory[32271] = 3'b110;
        rom_memory[32272] = 3'b110;
        rom_memory[32273] = 3'b110;
        rom_memory[32274] = 3'b110;
        rom_memory[32275] = 3'b110;
        rom_memory[32276] = 3'b110;
        rom_memory[32277] = 3'b110;
        rom_memory[32278] = 3'b110;
        rom_memory[32279] = 3'b110;
        rom_memory[32280] = 3'b110;
        rom_memory[32281] = 3'b110;
        rom_memory[32282] = 3'b110;
        rom_memory[32283] = 3'b110;
        rom_memory[32284] = 3'b110;
        rom_memory[32285] = 3'b110;
        rom_memory[32286] = 3'b110;
        rom_memory[32287] = 3'b110;
        rom_memory[32288] = 3'b110;
        rom_memory[32289] = 3'b110;
        rom_memory[32290] = 3'b110;
        rom_memory[32291] = 3'b111;
        rom_memory[32292] = 3'b110;
        rom_memory[32293] = 3'b000;
        rom_memory[32294] = 3'b000;
        rom_memory[32295] = 3'b000;
        rom_memory[32296] = 3'b000;
        rom_memory[32297] = 3'b000;
        rom_memory[32298] = 3'b000;
        rom_memory[32299] = 3'b000;
        rom_memory[32300] = 3'b000;
        rom_memory[32301] = 3'b100;
        rom_memory[32302] = 3'b110;
        rom_memory[32303] = 3'b110;
        rom_memory[32304] = 3'b100;
        rom_memory[32305] = 3'b000;
        rom_memory[32306] = 3'b100;
        rom_memory[32307] = 3'b110;
        rom_memory[32308] = 3'b111;
        rom_memory[32309] = 3'b110;
        rom_memory[32310] = 3'b110;
        rom_memory[32311] = 3'b110;
        rom_memory[32312] = 3'b110;
        rom_memory[32313] = 3'b110;
        rom_memory[32314] = 3'b110;
        rom_memory[32315] = 3'b110;
        rom_memory[32316] = 3'b110;
        rom_memory[32317] = 3'b110;
        rom_memory[32318] = 3'b110;
        rom_memory[32319] = 3'b110;
        rom_memory[32320] = 3'b110;
        rom_memory[32321] = 3'b110;
        rom_memory[32322] = 3'b110;
        rom_memory[32323] = 3'b110;
        rom_memory[32324] = 3'b110;
        rom_memory[32325] = 3'b110;
        rom_memory[32326] = 3'b110;
        rom_memory[32327] = 3'b110;
        rom_memory[32328] = 3'b110;
        rom_memory[32329] = 3'b110;
        rom_memory[32330] = 3'b110;
        rom_memory[32331] = 3'b110;
        rom_memory[32332] = 3'b110;
        rom_memory[32333] = 3'b110;
        rom_memory[32334] = 3'b110;
        rom_memory[32335] = 3'b110;
        rom_memory[32336] = 3'b110;
        rom_memory[32337] = 3'b110;
        rom_memory[32338] = 3'b110;
        rom_memory[32339] = 3'b110;
        rom_memory[32340] = 3'b110;
        rom_memory[32341] = 3'b110;
        rom_memory[32342] = 3'b110;
        rom_memory[32343] = 3'b110;
        rom_memory[32344] = 3'b111;
        rom_memory[32345] = 3'b111;
        rom_memory[32346] = 3'b111;
        rom_memory[32347] = 3'b111;
        rom_memory[32348] = 3'b111;
        rom_memory[32349] = 3'b111;
        rom_memory[32350] = 3'b111;
        rom_memory[32351] = 3'b111;
        rom_memory[32352] = 3'b111;
        rom_memory[32353] = 3'b111;
        rom_memory[32354] = 3'b111;
        rom_memory[32355] = 3'b111;
        rom_memory[32356] = 3'b111;
        rom_memory[32357] = 3'b111;
        rom_memory[32358] = 3'b111;
        rom_memory[32359] = 3'b111;
        rom_memory[32360] = 3'b111;
        rom_memory[32361] = 3'b111;
        rom_memory[32362] = 3'b111;
        rom_memory[32363] = 3'b111;
        rom_memory[32364] = 3'b111;
        rom_memory[32365] = 3'b111;
        rom_memory[32366] = 3'b111;
        rom_memory[32367] = 3'b111;
        rom_memory[32368] = 3'b111;
        rom_memory[32369] = 3'b111;
        rom_memory[32370] = 3'b111;
        rom_memory[32371] = 3'b111;
        rom_memory[32372] = 3'b111;
        rom_memory[32373] = 3'b111;
        rom_memory[32374] = 3'b111;
        rom_memory[32375] = 3'b111;
        rom_memory[32376] = 3'b111;
        rom_memory[32377] = 3'b111;
        rom_memory[32378] = 3'b111;
        rom_memory[32379] = 3'b111;
        rom_memory[32380] = 3'b111;
        rom_memory[32381] = 3'b111;
        rom_memory[32382] = 3'b111;
        rom_memory[32383] = 3'b111;
        rom_memory[32384] = 3'b111;
        rom_memory[32385] = 3'b111;
        rom_memory[32386] = 3'b111;
        rom_memory[32387] = 3'b111;
        rom_memory[32388] = 3'b111;
        rom_memory[32389] = 3'b111;
        rom_memory[32390] = 3'b111;
        rom_memory[32391] = 3'b111;
        rom_memory[32392] = 3'b111;
        rom_memory[32393] = 3'b111;
        rom_memory[32394] = 3'b111;
        rom_memory[32395] = 3'b111;
        rom_memory[32396] = 3'b111;
        rom_memory[32397] = 3'b111;
        rom_memory[32398] = 3'b111;
        rom_memory[32399] = 3'b111;
        rom_memory[32400] = 3'b110;
        rom_memory[32401] = 3'b110;
        rom_memory[32402] = 3'b110;
        rom_memory[32403] = 3'b110;
        rom_memory[32404] = 3'b110;
        rom_memory[32405] = 3'b110;
        rom_memory[32406] = 3'b110;
        rom_memory[32407] = 3'b110;
        rom_memory[32408] = 3'b111;
        rom_memory[32409] = 3'b111;
        rom_memory[32410] = 3'b111;
        rom_memory[32411] = 3'b111;
        rom_memory[32412] = 3'b111;
        rom_memory[32413] = 3'b111;
        rom_memory[32414] = 3'b111;
        rom_memory[32415] = 3'b111;
        rom_memory[32416] = 3'b111;
        rom_memory[32417] = 3'b111;
        rom_memory[32418] = 3'b111;
        rom_memory[32419] = 3'b111;
        rom_memory[32420] = 3'b110;
        rom_memory[32421] = 3'b110;
        rom_memory[32422] = 3'b110;
        rom_memory[32423] = 3'b110;
        rom_memory[32424] = 3'b110;
        rom_memory[32425] = 3'b110;
        rom_memory[32426] = 3'b111;
        rom_memory[32427] = 3'b111;
        rom_memory[32428] = 3'b111;
        rom_memory[32429] = 3'b111;
        rom_memory[32430] = 3'b111;
        rom_memory[32431] = 3'b111;
        rom_memory[32432] = 3'b111;
        rom_memory[32433] = 3'b111;
        rom_memory[32434] = 3'b111;
        rom_memory[32435] = 3'b111;
        rom_memory[32436] = 3'b111;
        rom_memory[32437] = 3'b111;
        rom_memory[32438] = 3'b111;
        rom_memory[32439] = 3'b110;
        rom_memory[32440] = 3'b111;
        rom_memory[32441] = 3'b110;
        rom_memory[32442] = 3'b110;
        rom_memory[32443] = 3'b110;
        rom_memory[32444] = 3'b110;
        rom_memory[32445] = 3'b111;
        rom_memory[32446] = 3'b111;
        rom_memory[32447] = 3'b111;
        rom_memory[32448] = 3'b111;
        rom_memory[32449] = 3'b111;
        rom_memory[32450] = 3'b111;
        rom_memory[32451] = 3'b111;
        rom_memory[32452] = 3'b111;
        rom_memory[32453] = 3'b111;
        rom_memory[32454] = 3'b111;
        rom_memory[32455] = 3'b111;
        rom_memory[32456] = 3'b111;
        rom_memory[32457] = 3'b111;
        rom_memory[32458] = 3'b111;
        rom_memory[32459] = 3'b111;
        rom_memory[32460] = 3'b111;
        rom_memory[32461] = 3'b111;
        rom_memory[32462] = 3'b000;
        rom_memory[32463] = 3'b000;
        rom_memory[32464] = 3'b000;
        rom_memory[32465] = 3'b000;
        rom_memory[32466] = 3'b000;
        rom_memory[32467] = 3'b000;
        rom_memory[32468] = 3'b000;
        rom_memory[32469] = 3'b000;
        rom_memory[32470] = 3'b000;
        rom_memory[32471] = 3'b000;
        rom_memory[32472] = 3'b000;
        rom_memory[32473] = 3'b111;
        rom_memory[32474] = 3'b111;
        rom_memory[32475] = 3'b111;
        rom_memory[32476] = 3'b111;
        rom_memory[32477] = 3'b111;
        rom_memory[32478] = 3'b110;
        rom_memory[32479] = 3'b110;
        rom_memory[32480] = 3'b110;
        rom_memory[32481] = 3'b111;
        rom_memory[32482] = 3'b110;
        rom_memory[32483] = 3'b100;
        rom_memory[32484] = 3'b110;
        rom_memory[32485] = 3'b110;
        rom_memory[32486] = 3'b111;
        rom_memory[32487] = 3'b111;
        rom_memory[32488] = 3'b111;
        rom_memory[32489] = 3'b110;
        rom_memory[32490] = 3'b000;
        rom_memory[32491] = 3'b000;
        rom_memory[32492] = 3'b110;
        rom_memory[32493] = 3'b111;
        rom_memory[32494] = 3'b111;
        rom_memory[32495] = 3'b100;
        rom_memory[32496] = 3'b110;
        rom_memory[32497] = 3'b111;
        rom_memory[32498] = 3'b111;
        rom_memory[32499] = 3'b110;
        rom_memory[32500] = 3'b110;
        rom_memory[32501] = 3'b110;
        rom_memory[32502] = 3'b110;
        rom_memory[32503] = 3'b110;
        rom_memory[32504] = 3'b110;
        rom_memory[32505] = 3'b110;
        rom_memory[32506] = 3'b110;
        rom_memory[32507] = 3'b110;
        rom_memory[32508] = 3'b110;
        rom_memory[32509] = 3'b110;
        rom_memory[32510] = 3'b110;
        rom_memory[32511] = 3'b110;
        rom_memory[32512] = 3'b110;
        rom_memory[32513] = 3'b110;
        rom_memory[32514] = 3'b110;
        rom_memory[32515] = 3'b110;
        rom_memory[32516] = 3'b110;
        rom_memory[32517] = 3'b110;
        rom_memory[32518] = 3'b110;
        rom_memory[32519] = 3'b110;
        rom_memory[32520] = 3'b110;
        rom_memory[32521] = 3'b110;
        rom_memory[32522] = 3'b110;
        rom_memory[32523] = 3'b110;
        rom_memory[32524] = 3'b110;
        rom_memory[32525] = 3'b110;
        rom_memory[32526] = 3'b110;
        rom_memory[32527] = 3'b110;
        rom_memory[32528] = 3'b110;
        rom_memory[32529] = 3'b110;
        rom_memory[32530] = 3'b110;
        rom_memory[32531] = 3'b110;
        rom_memory[32532] = 3'b110;
        rom_memory[32533] = 3'b110;
        rom_memory[32534] = 3'b000;
        rom_memory[32535] = 3'b000;
        rom_memory[32536] = 3'b000;
        rom_memory[32537] = 3'b000;
        rom_memory[32538] = 3'b000;
        rom_memory[32539] = 3'b000;
        rom_memory[32540] = 3'b100;
        rom_memory[32541] = 3'b100;
        rom_memory[32542] = 3'b100;
        rom_memory[32543] = 3'b100;
        rom_memory[32544] = 3'b110;
        rom_memory[32545] = 3'b100;
        rom_memory[32546] = 3'b000;
        rom_memory[32547] = 3'b100;
        rom_memory[32548] = 3'b110;
        rom_memory[32549] = 3'b111;
        rom_memory[32550] = 3'b110;
        rom_memory[32551] = 3'b110;
        rom_memory[32552] = 3'b110;
        rom_memory[32553] = 3'b110;
        rom_memory[32554] = 3'b110;
        rom_memory[32555] = 3'b110;
        rom_memory[32556] = 3'b110;
        rom_memory[32557] = 3'b110;
        rom_memory[32558] = 3'b110;
        rom_memory[32559] = 3'b110;
        rom_memory[32560] = 3'b110;
        rom_memory[32561] = 3'b110;
        rom_memory[32562] = 3'b110;
        rom_memory[32563] = 3'b110;
        rom_memory[32564] = 3'b110;
        rom_memory[32565] = 3'b110;
        rom_memory[32566] = 3'b110;
        rom_memory[32567] = 3'b110;
        rom_memory[32568] = 3'b110;
        rom_memory[32569] = 3'b110;
        rom_memory[32570] = 3'b110;
        rom_memory[32571] = 3'b110;
        rom_memory[32572] = 3'b110;
        rom_memory[32573] = 3'b110;
        rom_memory[32574] = 3'b110;
        rom_memory[32575] = 3'b110;
        rom_memory[32576] = 3'b110;
        rom_memory[32577] = 3'b110;
        rom_memory[32578] = 3'b110;
        rom_memory[32579] = 3'b110;
        rom_memory[32580] = 3'b110;
        rom_memory[32581] = 3'b110;
        rom_memory[32582] = 3'b110;
        rom_memory[32583] = 3'b110;
        rom_memory[32584] = 3'b111;
        rom_memory[32585] = 3'b111;
        rom_memory[32586] = 3'b111;
        rom_memory[32587] = 3'b111;
        rom_memory[32588] = 3'b111;
        rom_memory[32589] = 3'b111;
        rom_memory[32590] = 3'b111;
        rom_memory[32591] = 3'b111;
        rom_memory[32592] = 3'b111;
        rom_memory[32593] = 3'b111;
        rom_memory[32594] = 3'b111;
        rom_memory[32595] = 3'b111;
        rom_memory[32596] = 3'b111;
        rom_memory[32597] = 3'b111;
        rom_memory[32598] = 3'b111;
        rom_memory[32599] = 3'b111;
        rom_memory[32600] = 3'b111;
        rom_memory[32601] = 3'b111;
        rom_memory[32602] = 3'b111;
        rom_memory[32603] = 3'b111;
        rom_memory[32604] = 3'b111;
        rom_memory[32605] = 3'b111;
        rom_memory[32606] = 3'b111;
        rom_memory[32607] = 3'b111;
        rom_memory[32608] = 3'b111;
        rom_memory[32609] = 3'b111;
        rom_memory[32610] = 3'b111;
        rom_memory[32611] = 3'b111;
        rom_memory[32612] = 3'b111;
        rom_memory[32613] = 3'b111;
        rom_memory[32614] = 3'b111;
        rom_memory[32615] = 3'b111;
        rom_memory[32616] = 3'b111;
        rom_memory[32617] = 3'b111;
        rom_memory[32618] = 3'b111;
        rom_memory[32619] = 3'b111;
        rom_memory[32620] = 3'b111;
        rom_memory[32621] = 3'b111;
        rom_memory[32622] = 3'b111;
        rom_memory[32623] = 3'b111;
        rom_memory[32624] = 3'b111;
        rom_memory[32625] = 3'b111;
        rom_memory[32626] = 3'b111;
        rom_memory[32627] = 3'b111;
        rom_memory[32628] = 3'b111;
        rom_memory[32629] = 3'b111;
        rom_memory[32630] = 3'b111;
        rom_memory[32631] = 3'b111;
        rom_memory[32632] = 3'b111;
        rom_memory[32633] = 3'b111;
        rom_memory[32634] = 3'b111;
        rom_memory[32635] = 3'b111;
        rom_memory[32636] = 3'b111;
        rom_memory[32637] = 3'b111;
        rom_memory[32638] = 3'b111;
        rom_memory[32639] = 3'b111;
        rom_memory[32640] = 3'b110;
        rom_memory[32641] = 3'b110;
        rom_memory[32642] = 3'b110;
        rom_memory[32643] = 3'b110;
        rom_memory[32644] = 3'b110;
        rom_memory[32645] = 3'b110;
        rom_memory[32646] = 3'b110;
        rom_memory[32647] = 3'b111;
        rom_memory[32648] = 3'b111;
        rom_memory[32649] = 3'b111;
        rom_memory[32650] = 3'b111;
        rom_memory[32651] = 3'b111;
        rom_memory[32652] = 3'b111;
        rom_memory[32653] = 3'b111;
        rom_memory[32654] = 3'b111;
        rom_memory[32655] = 3'b111;
        rom_memory[32656] = 3'b111;
        rom_memory[32657] = 3'b111;
        rom_memory[32658] = 3'b111;
        rom_memory[32659] = 3'b111;
        rom_memory[32660] = 3'b110;
        rom_memory[32661] = 3'b110;
        rom_memory[32662] = 3'b110;
        rom_memory[32663] = 3'b110;
        rom_memory[32664] = 3'b110;
        rom_memory[32665] = 3'b110;
        rom_memory[32666] = 3'b111;
        rom_memory[32667] = 3'b111;
        rom_memory[32668] = 3'b111;
        rom_memory[32669] = 3'b111;
        rom_memory[32670] = 3'b111;
        rom_memory[32671] = 3'b111;
        rom_memory[32672] = 3'b111;
        rom_memory[32673] = 3'b111;
        rom_memory[32674] = 3'b111;
        rom_memory[32675] = 3'b111;
        rom_memory[32676] = 3'b110;
        rom_memory[32677] = 3'b110;
        rom_memory[32678] = 3'b110;
        rom_memory[32679] = 3'b110;
        rom_memory[32680] = 3'b110;
        rom_memory[32681] = 3'b110;
        rom_memory[32682] = 3'b110;
        rom_memory[32683] = 3'b110;
        rom_memory[32684] = 3'b110;
        rom_memory[32685] = 3'b111;
        rom_memory[32686] = 3'b111;
        rom_memory[32687] = 3'b111;
        rom_memory[32688] = 3'b111;
        rom_memory[32689] = 3'b111;
        rom_memory[32690] = 3'b111;
        rom_memory[32691] = 3'b111;
        rom_memory[32692] = 3'b111;
        rom_memory[32693] = 3'b111;
        rom_memory[32694] = 3'b111;
        rom_memory[32695] = 3'b111;
        rom_memory[32696] = 3'b111;
        rom_memory[32697] = 3'b111;
        rom_memory[32698] = 3'b111;
        rom_memory[32699] = 3'b111;
        rom_memory[32700] = 3'b111;
        rom_memory[32701] = 3'b111;
        rom_memory[32702] = 3'b000;
        rom_memory[32703] = 3'b000;
        rom_memory[32704] = 3'b000;
        rom_memory[32705] = 3'b000;
        rom_memory[32706] = 3'b000;
        rom_memory[32707] = 3'b000;
        rom_memory[32708] = 3'b000;
        rom_memory[32709] = 3'b000;
        rom_memory[32710] = 3'b000;
        rom_memory[32711] = 3'b000;
        rom_memory[32712] = 3'b111;
        rom_memory[32713] = 3'b111;
        rom_memory[32714] = 3'b111;
        rom_memory[32715] = 3'b111;
        rom_memory[32716] = 3'b111;
        rom_memory[32717] = 3'b111;
        rom_memory[32718] = 3'b111;
        rom_memory[32719] = 3'b111;
        rom_memory[32720] = 3'b111;
        rom_memory[32721] = 3'b111;
        rom_memory[32722] = 3'b111;
        rom_memory[32723] = 3'b110;
        rom_memory[32724] = 3'b110;
        rom_memory[32725] = 3'b100;
        rom_memory[32726] = 3'b111;
        rom_memory[32727] = 3'b111;
        rom_memory[32728] = 3'b110;
        rom_memory[32729] = 3'b000;
        rom_memory[32730] = 3'b000;
        rom_memory[32731] = 3'b000;
        rom_memory[32732] = 3'b111;
        rom_memory[32733] = 3'b111;
        rom_memory[32734] = 3'b111;
        rom_memory[32735] = 3'b111;
        rom_memory[32736] = 3'b111;
        rom_memory[32737] = 3'b111;
        rom_memory[32738] = 3'b111;
        rom_memory[32739] = 3'b110;
        rom_memory[32740] = 3'b110;
        rom_memory[32741] = 3'b110;
        rom_memory[32742] = 3'b110;
        rom_memory[32743] = 3'b110;
        rom_memory[32744] = 3'b110;
        rom_memory[32745] = 3'b110;
        rom_memory[32746] = 3'b110;
        rom_memory[32747] = 3'b110;
        rom_memory[32748] = 3'b110;
        rom_memory[32749] = 3'b110;
        rom_memory[32750] = 3'b110;
        rom_memory[32751] = 3'b110;
        rom_memory[32752] = 3'b110;
        rom_memory[32753] = 3'b110;
        rom_memory[32754] = 3'b110;
        rom_memory[32755] = 3'b110;
        rom_memory[32756] = 3'b110;
        rom_memory[32757] = 3'b110;
        rom_memory[32758] = 3'b110;
        rom_memory[32759] = 3'b110;
        rom_memory[32760] = 3'b110;
        rom_memory[32761] = 3'b110;
        rom_memory[32762] = 3'b110;
        rom_memory[32763] = 3'b110;
        rom_memory[32764] = 3'b110;
        rom_memory[32765] = 3'b110;
        rom_memory[32766] = 3'b110;
        rom_memory[32767] = 3'b110;
        rom_memory[32768] = 3'b110;
        rom_memory[32769] = 3'b110;
        rom_memory[32770] = 3'b110;
        rom_memory[32771] = 3'b110;
        rom_memory[32772] = 3'b110;
        rom_memory[32773] = 3'b110;
        rom_memory[32774] = 3'b110;
        rom_memory[32775] = 3'b000;
        rom_memory[32776] = 3'b000;
        rom_memory[32777] = 3'b000;
        rom_memory[32778] = 3'b000;
        rom_memory[32779] = 3'b000;
        rom_memory[32780] = 3'b000;
        rom_memory[32781] = 3'b110;
        rom_memory[32782] = 3'b100;
        rom_memory[32783] = 3'b000;
        rom_memory[32784] = 3'b100;
        rom_memory[32785] = 3'b110;
        rom_memory[32786] = 3'b100;
        rom_memory[32787] = 3'b000;
        rom_memory[32788] = 3'b100;
        rom_memory[32789] = 3'b100;
        rom_memory[32790] = 3'b111;
        rom_memory[32791] = 3'b110;
        rom_memory[32792] = 3'b110;
        rom_memory[32793] = 3'b110;
        rom_memory[32794] = 3'b110;
        rom_memory[32795] = 3'b110;
        rom_memory[32796] = 3'b110;
        rom_memory[32797] = 3'b110;
        rom_memory[32798] = 3'b110;
        rom_memory[32799] = 3'b110;
        rom_memory[32800] = 3'b110;
        rom_memory[32801] = 3'b110;
        rom_memory[32802] = 3'b110;
        rom_memory[32803] = 3'b110;
        rom_memory[32804] = 3'b110;
        rom_memory[32805] = 3'b110;
        rom_memory[32806] = 3'b110;
        rom_memory[32807] = 3'b110;
        rom_memory[32808] = 3'b110;
        rom_memory[32809] = 3'b110;
        rom_memory[32810] = 3'b110;
        rom_memory[32811] = 3'b110;
        rom_memory[32812] = 3'b110;
        rom_memory[32813] = 3'b110;
        rom_memory[32814] = 3'b110;
        rom_memory[32815] = 3'b110;
        rom_memory[32816] = 3'b110;
        rom_memory[32817] = 3'b110;
        rom_memory[32818] = 3'b110;
        rom_memory[32819] = 3'b110;
        rom_memory[32820] = 3'b110;
        rom_memory[32821] = 3'b110;
        rom_memory[32822] = 3'b110;
        rom_memory[32823] = 3'b110;
        rom_memory[32824] = 3'b111;
        rom_memory[32825] = 3'b111;
        rom_memory[32826] = 3'b111;
        rom_memory[32827] = 3'b111;
        rom_memory[32828] = 3'b111;
        rom_memory[32829] = 3'b111;
        rom_memory[32830] = 3'b111;
        rom_memory[32831] = 3'b111;
        rom_memory[32832] = 3'b111;
        rom_memory[32833] = 3'b111;
        rom_memory[32834] = 3'b111;
        rom_memory[32835] = 3'b111;
        rom_memory[32836] = 3'b111;
        rom_memory[32837] = 3'b111;
        rom_memory[32838] = 3'b111;
        rom_memory[32839] = 3'b111;
        rom_memory[32840] = 3'b111;
        rom_memory[32841] = 3'b111;
        rom_memory[32842] = 3'b111;
        rom_memory[32843] = 3'b111;
        rom_memory[32844] = 3'b111;
        rom_memory[32845] = 3'b111;
        rom_memory[32846] = 3'b111;
        rom_memory[32847] = 3'b111;
        rom_memory[32848] = 3'b111;
        rom_memory[32849] = 3'b111;
        rom_memory[32850] = 3'b111;
        rom_memory[32851] = 3'b111;
        rom_memory[32852] = 3'b111;
        rom_memory[32853] = 3'b111;
        rom_memory[32854] = 3'b111;
        rom_memory[32855] = 3'b111;
        rom_memory[32856] = 3'b111;
        rom_memory[32857] = 3'b111;
        rom_memory[32858] = 3'b111;
        rom_memory[32859] = 3'b111;
        rom_memory[32860] = 3'b111;
        rom_memory[32861] = 3'b111;
        rom_memory[32862] = 3'b111;
        rom_memory[32863] = 3'b111;
        rom_memory[32864] = 3'b111;
        rom_memory[32865] = 3'b111;
        rom_memory[32866] = 3'b111;
        rom_memory[32867] = 3'b111;
        rom_memory[32868] = 3'b111;
        rom_memory[32869] = 3'b111;
        rom_memory[32870] = 3'b111;
        rom_memory[32871] = 3'b111;
        rom_memory[32872] = 3'b111;
        rom_memory[32873] = 3'b111;
        rom_memory[32874] = 3'b111;
        rom_memory[32875] = 3'b111;
        rom_memory[32876] = 3'b111;
        rom_memory[32877] = 3'b111;
        rom_memory[32878] = 3'b111;
        rom_memory[32879] = 3'b111;
        rom_memory[32880] = 3'b110;
        rom_memory[32881] = 3'b110;
        rom_memory[32882] = 3'b110;
        rom_memory[32883] = 3'b110;
        rom_memory[32884] = 3'b110;
        rom_memory[32885] = 3'b110;
        rom_memory[32886] = 3'b110;
        rom_memory[32887] = 3'b111;
        rom_memory[32888] = 3'b111;
        rom_memory[32889] = 3'b111;
        rom_memory[32890] = 3'b111;
        rom_memory[32891] = 3'b111;
        rom_memory[32892] = 3'b111;
        rom_memory[32893] = 3'b111;
        rom_memory[32894] = 3'b111;
        rom_memory[32895] = 3'b111;
        rom_memory[32896] = 3'b111;
        rom_memory[32897] = 3'b111;
        rom_memory[32898] = 3'b111;
        rom_memory[32899] = 3'b111;
        rom_memory[32900] = 3'b110;
        rom_memory[32901] = 3'b110;
        rom_memory[32902] = 3'b110;
        rom_memory[32903] = 3'b110;
        rom_memory[32904] = 3'b110;
        rom_memory[32905] = 3'b111;
        rom_memory[32906] = 3'b111;
        rom_memory[32907] = 3'b111;
        rom_memory[32908] = 3'b111;
        rom_memory[32909] = 3'b111;
        rom_memory[32910] = 3'b111;
        rom_memory[32911] = 3'b111;
        rom_memory[32912] = 3'b111;
        rom_memory[32913] = 3'b111;
        rom_memory[32914] = 3'b111;
        rom_memory[32915] = 3'b110;
        rom_memory[32916] = 3'b110;
        rom_memory[32917] = 3'b110;
        rom_memory[32918] = 3'b110;
        rom_memory[32919] = 3'b110;
        rom_memory[32920] = 3'b110;
        rom_memory[32921] = 3'b110;
        rom_memory[32922] = 3'b110;
        rom_memory[32923] = 3'b110;
        rom_memory[32924] = 3'b110;
        rom_memory[32925] = 3'b110;
        rom_memory[32926] = 3'b111;
        rom_memory[32927] = 3'b111;
        rom_memory[32928] = 3'b111;
        rom_memory[32929] = 3'b111;
        rom_memory[32930] = 3'b111;
        rom_memory[32931] = 3'b111;
        rom_memory[32932] = 3'b111;
        rom_memory[32933] = 3'b111;
        rom_memory[32934] = 3'b111;
        rom_memory[32935] = 3'b111;
        rom_memory[32936] = 3'b111;
        rom_memory[32937] = 3'b111;
        rom_memory[32938] = 3'b111;
        rom_memory[32939] = 3'b111;
        rom_memory[32940] = 3'b111;
        rom_memory[32941] = 3'b111;
        rom_memory[32942] = 3'b000;
        rom_memory[32943] = 3'b000;
        rom_memory[32944] = 3'b000;
        rom_memory[32945] = 3'b000;
        rom_memory[32946] = 3'b000;
        rom_memory[32947] = 3'b000;
        rom_memory[32948] = 3'b000;
        rom_memory[32949] = 3'b000;
        rom_memory[32950] = 3'b000;
        rom_memory[32951] = 3'b111;
        rom_memory[32952] = 3'b111;
        rom_memory[32953] = 3'b111;
        rom_memory[32954] = 3'b111;
        rom_memory[32955] = 3'b110;
        rom_memory[32956] = 3'b111;
        rom_memory[32957] = 3'b111;
        rom_memory[32958] = 3'b111;
        rom_memory[32959] = 3'b111;
        rom_memory[32960] = 3'b111;
        rom_memory[32961] = 3'b110;
        rom_memory[32962] = 3'b110;
        rom_memory[32963] = 3'b100;
        rom_memory[32964] = 3'b100;
        rom_memory[32965] = 3'b110;
        rom_memory[32966] = 3'b110;
        rom_memory[32967] = 3'b110;
        rom_memory[32968] = 3'b100;
        rom_memory[32969] = 3'b100;
        rom_memory[32970] = 3'b110;
        rom_memory[32971] = 3'b100;
        rom_memory[32972] = 3'b111;
        rom_memory[32973] = 3'b111;
        rom_memory[32974] = 3'b111;
        rom_memory[32975] = 3'b111;
        rom_memory[32976] = 3'b111;
        rom_memory[32977] = 3'b110;
        rom_memory[32978] = 3'b110;
        rom_memory[32979] = 3'b110;
        rom_memory[32980] = 3'b110;
        rom_memory[32981] = 3'b110;
        rom_memory[32982] = 3'b110;
        rom_memory[32983] = 3'b110;
        rom_memory[32984] = 3'b110;
        rom_memory[32985] = 3'b110;
        rom_memory[32986] = 3'b110;
        rom_memory[32987] = 3'b110;
        rom_memory[32988] = 3'b110;
        rom_memory[32989] = 3'b110;
        rom_memory[32990] = 3'b110;
        rom_memory[32991] = 3'b110;
        rom_memory[32992] = 3'b110;
        rom_memory[32993] = 3'b110;
        rom_memory[32994] = 3'b110;
        rom_memory[32995] = 3'b110;
        rom_memory[32996] = 3'b110;
        rom_memory[32997] = 3'b110;
        rom_memory[32998] = 3'b110;
        rom_memory[32999] = 3'b110;
        rom_memory[33000] = 3'b110;
        rom_memory[33001] = 3'b110;
        rom_memory[33002] = 3'b110;
        rom_memory[33003] = 3'b110;
        rom_memory[33004] = 3'b110;
        rom_memory[33005] = 3'b110;
        rom_memory[33006] = 3'b110;
        rom_memory[33007] = 3'b110;
        rom_memory[33008] = 3'b110;
        rom_memory[33009] = 3'b110;
        rom_memory[33010] = 3'b110;
        rom_memory[33011] = 3'b110;
        rom_memory[33012] = 3'b110;
        rom_memory[33013] = 3'b110;
        rom_memory[33014] = 3'b110;
        rom_memory[33015] = 3'b110;
        rom_memory[33016] = 3'b000;
        rom_memory[33017] = 3'b000;
        rom_memory[33018] = 3'b000;
        rom_memory[33019] = 3'b000;
        rom_memory[33020] = 3'b000;
        rom_memory[33021] = 3'b000;
        rom_memory[33022] = 3'b110;
        rom_memory[33023] = 3'b100;
        rom_memory[33024] = 3'b000;
        rom_memory[33025] = 3'b100;
        rom_memory[33026] = 3'b110;
        rom_memory[33027] = 3'b100;
        rom_memory[33028] = 3'b000;
        rom_memory[33029] = 3'b000;
        rom_memory[33030] = 3'b100;
        rom_memory[33031] = 3'b111;
        rom_memory[33032] = 3'b110;
        rom_memory[33033] = 3'b110;
        rom_memory[33034] = 3'b110;
        rom_memory[33035] = 3'b110;
        rom_memory[33036] = 3'b110;
        rom_memory[33037] = 3'b110;
        rom_memory[33038] = 3'b110;
        rom_memory[33039] = 3'b110;
        rom_memory[33040] = 3'b110;
        rom_memory[33041] = 3'b110;
        rom_memory[33042] = 3'b110;
        rom_memory[33043] = 3'b110;
        rom_memory[33044] = 3'b110;
        rom_memory[33045] = 3'b110;
        rom_memory[33046] = 3'b110;
        rom_memory[33047] = 3'b110;
        rom_memory[33048] = 3'b110;
        rom_memory[33049] = 3'b110;
        rom_memory[33050] = 3'b110;
        rom_memory[33051] = 3'b110;
        rom_memory[33052] = 3'b110;
        rom_memory[33053] = 3'b110;
        rom_memory[33054] = 3'b110;
        rom_memory[33055] = 3'b110;
        rom_memory[33056] = 3'b110;
        rom_memory[33057] = 3'b110;
        rom_memory[33058] = 3'b110;
        rom_memory[33059] = 3'b110;
        rom_memory[33060] = 3'b110;
        rom_memory[33061] = 3'b110;
        rom_memory[33062] = 3'b110;
        rom_memory[33063] = 3'b110;
        rom_memory[33064] = 3'b110;
        rom_memory[33065] = 3'b110;
        rom_memory[33066] = 3'b111;
        rom_memory[33067] = 3'b111;
        rom_memory[33068] = 3'b111;
        rom_memory[33069] = 3'b111;
        rom_memory[33070] = 3'b111;
        rom_memory[33071] = 3'b111;
        rom_memory[33072] = 3'b111;
        rom_memory[33073] = 3'b111;
        rom_memory[33074] = 3'b111;
        rom_memory[33075] = 3'b111;
        rom_memory[33076] = 3'b111;
        rom_memory[33077] = 3'b111;
        rom_memory[33078] = 3'b111;
        rom_memory[33079] = 3'b111;
        rom_memory[33080] = 3'b111;
        rom_memory[33081] = 3'b111;
        rom_memory[33082] = 3'b111;
        rom_memory[33083] = 3'b111;
        rom_memory[33084] = 3'b111;
        rom_memory[33085] = 3'b111;
        rom_memory[33086] = 3'b111;
        rom_memory[33087] = 3'b111;
        rom_memory[33088] = 3'b111;
        rom_memory[33089] = 3'b111;
        rom_memory[33090] = 3'b111;
        rom_memory[33091] = 3'b111;
        rom_memory[33092] = 3'b111;
        rom_memory[33093] = 3'b111;
        rom_memory[33094] = 3'b111;
        rom_memory[33095] = 3'b111;
        rom_memory[33096] = 3'b111;
        rom_memory[33097] = 3'b111;
        rom_memory[33098] = 3'b111;
        rom_memory[33099] = 3'b111;
        rom_memory[33100] = 3'b111;
        rom_memory[33101] = 3'b111;
        rom_memory[33102] = 3'b111;
        rom_memory[33103] = 3'b111;
        rom_memory[33104] = 3'b111;
        rom_memory[33105] = 3'b111;
        rom_memory[33106] = 3'b111;
        rom_memory[33107] = 3'b111;
        rom_memory[33108] = 3'b111;
        rom_memory[33109] = 3'b111;
        rom_memory[33110] = 3'b111;
        rom_memory[33111] = 3'b111;
        rom_memory[33112] = 3'b111;
        rom_memory[33113] = 3'b111;
        rom_memory[33114] = 3'b111;
        rom_memory[33115] = 3'b111;
        rom_memory[33116] = 3'b111;
        rom_memory[33117] = 3'b111;
        rom_memory[33118] = 3'b111;
        rom_memory[33119] = 3'b111;
        rom_memory[33120] = 3'b110;
        rom_memory[33121] = 3'b110;
        rom_memory[33122] = 3'b110;
        rom_memory[33123] = 3'b110;
        rom_memory[33124] = 3'b110;
        rom_memory[33125] = 3'b110;
        rom_memory[33126] = 3'b111;
        rom_memory[33127] = 3'b111;
        rom_memory[33128] = 3'b111;
        rom_memory[33129] = 3'b111;
        rom_memory[33130] = 3'b111;
        rom_memory[33131] = 3'b111;
        rom_memory[33132] = 3'b111;
        rom_memory[33133] = 3'b111;
        rom_memory[33134] = 3'b111;
        rom_memory[33135] = 3'b111;
        rom_memory[33136] = 3'b111;
        rom_memory[33137] = 3'b111;
        rom_memory[33138] = 3'b111;
        rom_memory[33139] = 3'b111;
        rom_memory[33140] = 3'b110;
        rom_memory[33141] = 3'b110;
        rom_memory[33142] = 3'b110;
        rom_memory[33143] = 3'b110;
        rom_memory[33144] = 3'b110;
        rom_memory[33145] = 3'b110;
        rom_memory[33146] = 3'b111;
        rom_memory[33147] = 3'b111;
        rom_memory[33148] = 3'b111;
        rom_memory[33149] = 3'b111;
        rom_memory[33150] = 3'b111;
        rom_memory[33151] = 3'b111;
        rom_memory[33152] = 3'b111;
        rom_memory[33153] = 3'b111;
        rom_memory[33154] = 3'b111;
        rom_memory[33155] = 3'b110;
        rom_memory[33156] = 3'b110;
        rom_memory[33157] = 3'b110;
        rom_memory[33158] = 3'b110;
        rom_memory[33159] = 3'b110;
        rom_memory[33160] = 3'b110;
        rom_memory[33161] = 3'b110;
        rom_memory[33162] = 3'b110;
        rom_memory[33163] = 3'b110;
        rom_memory[33164] = 3'b110;
        rom_memory[33165] = 3'b110;
        rom_memory[33166] = 3'b111;
        rom_memory[33167] = 3'b111;
        rom_memory[33168] = 3'b111;
        rom_memory[33169] = 3'b111;
        rom_memory[33170] = 3'b111;
        rom_memory[33171] = 3'b111;
        rom_memory[33172] = 3'b111;
        rom_memory[33173] = 3'b111;
        rom_memory[33174] = 3'b111;
        rom_memory[33175] = 3'b111;
        rom_memory[33176] = 3'b111;
        rom_memory[33177] = 3'b111;
        rom_memory[33178] = 3'b111;
        rom_memory[33179] = 3'b111;
        rom_memory[33180] = 3'b111;
        rom_memory[33181] = 3'b111;
        rom_memory[33182] = 3'b000;
        rom_memory[33183] = 3'b000;
        rom_memory[33184] = 3'b000;
        rom_memory[33185] = 3'b000;
        rom_memory[33186] = 3'b000;
        rom_memory[33187] = 3'b000;
        rom_memory[33188] = 3'b000;
        rom_memory[33189] = 3'b000;
        rom_memory[33190] = 3'b000;
        rom_memory[33191] = 3'b000;
        rom_memory[33192] = 3'b110;
        rom_memory[33193] = 3'b110;
        rom_memory[33194] = 3'b111;
        rom_memory[33195] = 3'b111;
        rom_memory[33196] = 3'b111;
        rom_memory[33197] = 3'b111;
        rom_memory[33198] = 3'b111;
        rom_memory[33199] = 3'b111;
        rom_memory[33200] = 3'b110;
        rom_memory[33201] = 3'b000;
        rom_memory[33202] = 3'b000;
        rom_memory[33203] = 3'b000;
        rom_memory[33204] = 3'b000;
        rom_memory[33205] = 3'b100;
        rom_memory[33206] = 3'b111;
        rom_memory[33207] = 3'b111;
        rom_memory[33208] = 3'b000;
        rom_memory[33209] = 3'b000;
        rom_memory[33210] = 3'b100;
        rom_memory[33211] = 3'b111;
        rom_memory[33212] = 3'b111;
        rom_memory[33213] = 3'b111;
        rom_memory[33214] = 3'b111;
        rom_memory[33215] = 3'b111;
        rom_memory[33216] = 3'b111;
        rom_memory[33217] = 3'b111;
        rom_memory[33218] = 3'b110;
        rom_memory[33219] = 3'b110;
        rom_memory[33220] = 3'b110;
        rom_memory[33221] = 3'b110;
        rom_memory[33222] = 3'b110;
        rom_memory[33223] = 3'b110;
        rom_memory[33224] = 3'b110;
        rom_memory[33225] = 3'b110;
        rom_memory[33226] = 3'b110;
        rom_memory[33227] = 3'b110;
        rom_memory[33228] = 3'b110;
        rom_memory[33229] = 3'b110;
        rom_memory[33230] = 3'b110;
        rom_memory[33231] = 3'b110;
        rom_memory[33232] = 3'b110;
        rom_memory[33233] = 3'b110;
        rom_memory[33234] = 3'b110;
        rom_memory[33235] = 3'b110;
        rom_memory[33236] = 3'b110;
        rom_memory[33237] = 3'b110;
        rom_memory[33238] = 3'b110;
        rom_memory[33239] = 3'b110;
        rom_memory[33240] = 3'b110;
        rom_memory[33241] = 3'b110;
        rom_memory[33242] = 3'b110;
        rom_memory[33243] = 3'b110;
        rom_memory[33244] = 3'b110;
        rom_memory[33245] = 3'b110;
        rom_memory[33246] = 3'b110;
        rom_memory[33247] = 3'b110;
        rom_memory[33248] = 3'b110;
        rom_memory[33249] = 3'b110;
        rom_memory[33250] = 3'b110;
        rom_memory[33251] = 3'b110;
        rom_memory[33252] = 3'b110;
        rom_memory[33253] = 3'b110;
        rom_memory[33254] = 3'b110;
        rom_memory[33255] = 3'b110;
        rom_memory[33256] = 3'b110;
        rom_memory[33257] = 3'b000;
        rom_memory[33258] = 3'b000;
        rom_memory[33259] = 3'b000;
        rom_memory[33260] = 3'b000;
        rom_memory[33261] = 3'b000;
        rom_memory[33262] = 3'b000;
        rom_memory[33263] = 3'b110;
        rom_memory[33264] = 3'b100;
        rom_memory[33265] = 3'b000;
        rom_memory[33266] = 3'b100;
        rom_memory[33267] = 3'b110;
        rom_memory[33268] = 3'b100;
        rom_memory[33269] = 3'b000;
        rom_memory[33270] = 3'b000;
        rom_memory[33271] = 3'b110;
        rom_memory[33272] = 3'b110;
        rom_memory[33273] = 3'b110;
        rom_memory[33274] = 3'b110;
        rom_memory[33275] = 3'b110;
        rom_memory[33276] = 3'b110;
        rom_memory[33277] = 3'b110;
        rom_memory[33278] = 3'b110;
        rom_memory[33279] = 3'b110;
        rom_memory[33280] = 3'b110;
        rom_memory[33281] = 3'b110;
        rom_memory[33282] = 3'b110;
        rom_memory[33283] = 3'b110;
        rom_memory[33284] = 3'b110;
        rom_memory[33285] = 3'b110;
        rom_memory[33286] = 3'b110;
        rom_memory[33287] = 3'b110;
        rom_memory[33288] = 3'b110;
        rom_memory[33289] = 3'b110;
        rom_memory[33290] = 3'b110;
        rom_memory[33291] = 3'b110;
        rom_memory[33292] = 3'b110;
        rom_memory[33293] = 3'b110;
        rom_memory[33294] = 3'b110;
        rom_memory[33295] = 3'b110;
        rom_memory[33296] = 3'b110;
        rom_memory[33297] = 3'b110;
        rom_memory[33298] = 3'b110;
        rom_memory[33299] = 3'b110;
        rom_memory[33300] = 3'b110;
        rom_memory[33301] = 3'b110;
        rom_memory[33302] = 3'b110;
        rom_memory[33303] = 3'b110;
        rom_memory[33304] = 3'b110;
        rom_memory[33305] = 3'b110;
        rom_memory[33306] = 3'b111;
        rom_memory[33307] = 3'b111;
        rom_memory[33308] = 3'b111;
        rom_memory[33309] = 3'b111;
        rom_memory[33310] = 3'b111;
        rom_memory[33311] = 3'b111;
        rom_memory[33312] = 3'b111;
        rom_memory[33313] = 3'b111;
        rom_memory[33314] = 3'b111;
        rom_memory[33315] = 3'b111;
        rom_memory[33316] = 3'b111;
        rom_memory[33317] = 3'b111;
        rom_memory[33318] = 3'b111;
        rom_memory[33319] = 3'b111;
        rom_memory[33320] = 3'b111;
        rom_memory[33321] = 3'b111;
        rom_memory[33322] = 3'b111;
        rom_memory[33323] = 3'b111;
        rom_memory[33324] = 3'b111;
        rom_memory[33325] = 3'b111;
        rom_memory[33326] = 3'b111;
        rom_memory[33327] = 3'b111;
        rom_memory[33328] = 3'b111;
        rom_memory[33329] = 3'b111;
        rom_memory[33330] = 3'b111;
        rom_memory[33331] = 3'b111;
        rom_memory[33332] = 3'b111;
        rom_memory[33333] = 3'b111;
        rom_memory[33334] = 3'b111;
        rom_memory[33335] = 3'b111;
        rom_memory[33336] = 3'b111;
        rom_memory[33337] = 3'b111;
        rom_memory[33338] = 3'b111;
        rom_memory[33339] = 3'b111;
        rom_memory[33340] = 3'b111;
        rom_memory[33341] = 3'b111;
        rom_memory[33342] = 3'b111;
        rom_memory[33343] = 3'b111;
        rom_memory[33344] = 3'b111;
        rom_memory[33345] = 3'b111;
        rom_memory[33346] = 3'b111;
        rom_memory[33347] = 3'b111;
        rom_memory[33348] = 3'b111;
        rom_memory[33349] = 3'b111;
        rom_memory[33350] = 3'b111;
        rom_memory[33351] = 3'b111;
        rom_memory[33352] = 3'b111;
        rom_memory[33353] = 3'b111;
        rom_memory[33354] = 3'b111;
        rom_memory[33355] = 3'b111;
        rom_memory[33356] = 3'b111;
        rom_memory[33357] = 3'b111;
        rom_memory[33358] = 3'b111;
        rom_memory[33359] = 3'b111;
        rom_memory[33360] = 3'b110;
        rom_memory[33361] = 3'b110;
        rom_memory[33362] = 3'b110;
        rom_memory[33363] = 3'b110;
        rom_memory[33364] = 3'b110;
        rom_memory[33365] = 3'b110;
        rom_memory[33366] = 3'b111;
        rom_memory[33367] = 3'b111;
        rom_memory[33368] = 3'b111;
        rom_memory[33369] = 3'b111;
        rom_memory[33370] = 3'b111;
        rom_memory[33371] = 3'b111;
        rom_memory[33372] = 3'b111;
        rom_memory[33373] = 3'b111;
        rom_memory[33374] = 3'b111;
        rom_memory[33375] = 3'b111;
        rom_memory[33376] = 3'b111;
        rom_memory[33377] = 3'b111;
        rom_memory[33378] = 3'b111;
        rom_memory[33379] = 3'b111;
        rom_memory[33380] = 3'b111;
        rom_memory[33381] = 3'b110;
        rom_memory[33382] = 3'b110;
        rom_memory[33383] = 3'b110;
        rom_memory[33384] = 3'b110;
        rom_memory[33385] = 3'b110;
        rom_memory[33386] = 3'b111;
        rom_memory[33387] = 3'b111;
        rom_memory[33388] = 3'b111;
        rom_memory[33389] = 3'b111;
        rom_memory[33390] = 3'b111;
        rom_memory[33391] = 3'b111;
        rom_memory[33392] = 3'b111;
        rom_memory[33393] = 3'b111;
        rom_memory[33394] = 3'b111;
        rom_memory[33395] = 3'b110;
        rom_memory[33396] = 3'b110;
        rom_memory[33397] = 3'b110;
        rom_memory[33398] = 3'b110;
        rom_memory[33399] = 3'b110;
        rom_memory[33400] = 3'b110;
        rom_memory[33401] = 3'b110;
        rom_memory[33402] = 3'b110;
        rom_memory[33403] = 3'b110;
        rom_memory[33404] = 3'b110;
        rom_memory[33405] = 3'b110;
        rom_memory[33406] = 3'b110;
        rom_memory[33407] = 3'b111;
        rom_memory[33408] = 3'b111;
        rom_memory[33409] = 3'b111;
        rom_memory[33410] = 3'b111;
        rom_memory[33411] = 3'b111;
        rom_memory[33412] = 3'b111;
        rom_memory[33413] = 3'b111;
        rom_memory[33414] = 3'b111;
        rom_memory[33415] = 3'b111;
        rom_memory[33416] = 3'b111;
        rom_memory[33417] = 3'b111;
        rom_memory[33418] = 3'b111;
        rom_memory[33419] = 3'b111;
        rom_memory[33420] = 3'b111;
        rom_memory[33421] = 3'b111;
        rom_memory[33422] = 3'b000;
        rom_memory[33423] = 3'b000;
        rom_memory[33424] = 3'b000;
        rom_memory[33425] = 3'b000;
        rom_memory[33426] = 3'b000;
        rom_memory[33427] = 3'b000;
        rom_memory[33428] = 3'b000;
        rom_memory[33429] = 3'b000;
        rom_memory[33430] = 3'b000;
        rom_memory[33431] = 3'b110;
        rom_memory[33432] = 3'b110;
        rom_memory[33433] = 3'b110;
        rom_memory[33434] = 3'b110;
        rom_memory[33435] = 3'b110;
        rom_memory[33436] = 3'b111;
        rom_memory[33437] = 3'b111;
        rom_memory[33438] = 3'b111;
        rom_memory[33439] = 3'b000;
        rom_memory[33440] = 3'b000;
        rom_memory[33441] = 3'b000;
        rom_memory[33442] = 3'b000;
        rom_memory[33443] = 3'b000;
        rom_memory[33444] = 3'b000;
        rom_memory[33445] = 3'b000;
        rom_memory[33446] = 3'b111;
        rom_memory[33447] = 3'b111;
        rom_memory[33448] = 3'b000;
        rom_memory[33449] = 3'b000;
        rom_memory[33450] = 3'b000;
        rom_memory[33451] = 3'b100;
        rom_memory[33452] = 3'b100;
        rom_memory[33453] = 3'b111;
        rom_memory[33454] = 3'b111;
        rom_memory[33455] = 3'b111;
        rom_memory[33456] = 3'b111;
        rom_memory[33457] = 3'b111;
        rom_memory[33458] = 3'b111;
        rom_memory[33459] = 3'b110;
        rom_memory[33460] = 3'b110;
        rom_memory[33461] = 3'b110;
        rom_memory[33462] = 3'b110;
        rom_memory[33463] = 3'b110;
        rom_memory[33464] = 3'b110;
        rom_memory[33465] = 3'b110;
        rom_memory[33466] = 3'b110;
        rom_memory[33467] = 3'b110;
        rom_memory[33468] = 3'b110;
        rom_memory[33469] = 3'b110;
        rom_memory[33470] = 3'b110;
        rom_memory[33471] = 3'b110;
        rom_memory[33472] = 3'b110;
        rom_memory[33473] = 3'b110;
        rom_memory[33474] = 3'b110;
        rom_memory[33475] = 3'b110;
        rom_memory[33476] = 3'b110;
        rom_memory[33477] = 3'b110;
        rom_memory[33478] = 3'b110;
        rom_memory[33479] = 3'b110;
        rom_memory[33480] = 3'b110;
        rom_memory[33481] = 3'b110;
        rom_memory[33482] = 3'b110;
        rom_memory[33483] = 3'b110;
        rom_memory[33484] = 3'b110;
        rom_memory[33485] = 3'b110;
        rom_memory[33486] = 3'b110;
        rom_memory[33487] = 3'b110;
        rom_memory[33488] = 3'b110;
        rom_memory[33489] = 3'b110;
        rom_memory[33490] = 3'b110;
        rom_memory[33491] = 3'b110;
        rom_memory[33492] = 3'b110;
        rom_memory[33493] = 3'b110;
        rom_memory[33494] = 3'b110;
        rom_memory[33495] = 3'b110;
        rom_memory[33496] = 3'b110;
        rom_memory[33497] = 3'b110;
        rom_memory[33498] = 3'b000;
        rom_memory[33499] = 3'b000;
        rom_memory[33500] = 3'b000;
        rom_memory[33501] = 3'b000;
        rom_memory[33502] = 3'b000;
        rom_memory[33503] = 3'b000;
        rom_memory[33504] = 3'b110;
        rom_memory[33505] = 3'b100;
        rom_memory[33506] = 3'b000;
        rom_memory[33507] = 3'b100;
        rom_memory[33508] = 3'b110;
        rom_memory[33509] = 3'b100;
        rom_memory[33510] = 3'b000;
        rom_memory[33511] = 3'b100;
        rom_memory[33512] = 3'b100;
        rom_memory[33513] = 3'b111;
        rom_memory[33514] = 3'b110;
        rom_memory[33515] = 3'b110;
        rom_memory[33516] = 3'b110;
        rom_memory[33517] = 3'b110;
        rom_memory[33518] = 3'b110;
        rom_memory[33519] = 3'b110;
        rom_memory[33520] = 3'b110;
        rom_memory[33521] = 3'b110;
        rom_memory[33522] = 3'b110;
        rom_memory[33523] = 3'b110;
        rom_memory[33524] = 3'b110;
        rom_memory[33525] = 3'b110;
        rom_memory[33526] = 3'b110;
        rom_memory[33527] = 3'b110;
        rom_memory[33528] = 3'b110;
        rom_memory[33529] = 3'b110;
        rom_memory[33530] = 3'b110;
        rom_memory[33531] = 3'b110;
        rom_memory[33532] = 3'b110;
        rom_memory[33533] = 3'b110;
        rom_memory[33534] = 3'b110;
        rom_memory[33535] = 3'b110;
        rom_memory[33536] = 3'b110;
        rom_memory[33537] = 3'b110;
        rom_memory[33538] = 3'b110;
        rom_memory[33539] = 3'b110;
        rom_memory[33540] = 3'b110;
        rom_memory[33541] = 3'b110;
        rom_memory[33542] = 3'b110;
        rom_memory[33543] = 3'b110;
        rom_memory[33544] = 3'b110;
        rom_memory[33545] = 3'b110;
        rom_memory[33546] = 3'b111;
        rom_memory[33547] = 3'b111;
        rom_memory[33548] = 3'b111;
        rom_memory[33549] = 3'b111;
        rom_memory[33550] = 3'b111;
        rom_memory[33551] = 3'b111;
        rom_memory[33552] = 3'b111;
        rom_memory[33553] = 3'b111;
        rom_memory[33554] = 3'b111;
        rom_memory[33555] = 3'b111;
        rom_memory[33556] = 3'b111;
        rom_memory[33557] = 3'b111;
        rom_memory[33558] = 3'b111;
        rom_memory[33559] = 3'b111;
        rom_memory[33560] = 3'b111;
        rom_memory[33561] = 3'b111;
        rom_memory[33562] = 3'b111;
        rom_memory[33563] = 3'b111;
        rom_memory[33564] = 3'b111;
        rom_memory[33565] = 3'b111;
        rom_memory[33566] = 3'b111;
        rom_memory[33567] = 3'b111;
        rom_memory[33568] = 3'b111;
        rom_memory[33569] = 3'b111;
        rom_memory[33570] = 3'b111;
        rom_memory[33571] = 3'b111;
        rom_memory[33572] = 3'b111;
        rom_memory[33573] = 3'b111;
        rom_memory[33574] = 3'b111;
        rom_memory[33575] = 3'b111;
        rom_memory[33576] = 3'b111;
        rom_memory[33577] = 3'b111;
        rom_memory[33578] = 3'b111;
        rom_memory[33579] = 3'b111;
        rom_memory[33580] = 3'b111;
        rom_memory[33581] = 3'b111;
        rom_memory[33582] = 3'b111;
        rom_memory[33583] = 3'b111;
        rom_memory[33584] = 3'b111;
        rom_memory[33585] = 3'b111;
        rom_memory[33586] = 3'b111;
        rom_memory[33587] = 3'b111;
        rom_memory[33588] = 3'b111;
        rom_memory[33589] = 3'b111;
        rom_memory[33590] = 3'b111;
        rom_memory[33591] = 3'b111;
        rom_memory[33592] = 3'b111;
        rom_memory[33593] = 3'b111;
        rom_memory[33594] = 3'b111;
        rom_memory[33595] = 3'b111;
        rom_memory[33596] = 3'b111;
        rom_memory[33597] = 3'b111;
        rom_memory[33598] = 3'b111;
        rom_memory[33599] = 3'b111;
        rom_memory[33600] = 3'b110;
        rom_memory[33601] = 3'b110;
        rom_memory[33602] = 3'b110;
        rom_memory[33603] = 3'b110;
        rom_memory[33604] = 3'b110;
        rom_memory[33605] = 3'b110;
        rom_memory[33606] = 3'b111;
        rom_memory[33607] = 3'b111;
        rom_memory[33608] = 3'b111;
        rom_memory[33609] = 3'b111;
        rom_memory[33610] = 3'b111;
        rom_memory[33611] = 3'b111;
        rom_memory[33612] = 3'b111;
        rom_memory[33613] = 3'b111;
        rom_memory[33614] = 3'b111;
        rom_memory[33615] = 3'b111;
        rom_memory[33616] = 3'b111;
        rom_memory[33617] = 3'b111;
        rom_memory[33618] = 3'b111;
        rom_memory[33619] = 3'b111;
        rom_memory[33620] = 3'b111;
        rom_memory[33621] = 3'b110;
        rom_memory[33622] = 3'b110;
        rom_memory[33623] = 3'b110;
        rom_memory[33624] = 3'b111;
        rom_memory[33625] = 3'b110;
        rom_memory[33626] = 3'b111;
        rom_memory[33627] = 3'b111;
        rom_memory[33628] = 3'b111;
        rom_memory[33629] = 3'b111;
        rom_memory[33630] = 3'b111;
        rom_memory[33631] = 3'b111;
        rom_memory[33632] = 3'b111;
        rom_memory[33633] = 3'b111;
        rom_memory[33634] = 3'b110;
        rom_memory[33635] = 3'b110;
        rom_memory[33636] = 3'b110;
        rom_memory[33637] = 3'b110;
        rom_memory[33638] = 3'b110;
        rom_memory[33639] = 3'b110;
        rom_memory[33640] = 3'b110;
        rom_memory[33641] = 3'b110;
        rom_memory[33642] = 3'b110;
        rom_memory[33643] = 3'b110;
        rom_memory[33644] = 3'b110;
        rom_memory[33645] = 3'b110;
        rom_memory[33646] = 3'b111;
        rom_memory[33647] = 3'b111;
        rom_memory[33648] = 3'b111;
        rom_memory[33649] = 3'b111;
        rom_memory[33650] = 3'b111;
        rom_memory[33651] = 3'b111;
        rom_memory[33652] = 3'b111;
        rom_memory[33653] = 3'b111;
        rom_memory[33654] = 3'b111;
        rom_memory[33655] = 3'b111;
        rom_memory[33656] = 3'b111;
        rom_memory[33657] = 3'b111;
        rom_memory[33658] = 3'b111;
        rom_memory[33659] = 3'b111;
        rom_memory[33660] = 3'b111;
        rom_memory[33661] = 3'b111;
        rom_memory[33662] = 3'b000;
        rom_memory[33663] = 3'b000;
        rom_memory[33664] = 3'b000;
        rom_memory[33665] = 3'b000;
        rom_memory[33666] = 3'b000;
        rom_memory[33667] = 3'b000;
        rom_memory[33668] = 3'b000;
        rom_memory[33669] = 3'b000;
        rom_memory[33670] = 3'b111;
        rom_memory[33671] = 3'b110;
        rom_memory[33672] = 3'b110;
        rom_memory[33673] = 3'b110;
        rom_memory[33674] = 3'b110;
        rom_memory[33675] = 3'b100;
        rom_memory[33676] = 3'b110;
        rom_memory[33677] = 3'b111;
        rom_memory[33678] = 3'b111;
        rom_memory[33679] = 3'b000;
        rom_memory[33680] = 3'b000;
        rom_memory[33681] = 3'b000;
        rom_memory[33682] = 3'b000;
        rom_memory[33683] = 3'b000;
        rom_memory[33684] = 3'b000;
        rom_memory[33685] = 3'b000;
        rom_memory[33686] = 3'b000;
        rom_memory[33687] = 3'b110;
        rom_memory[33688] = 3'b100;
        rom_memory[33689] = 3'b100;
        rom_memory[33690] = 3'b100;
        rom_memory[33691] = 3'b110;
        rom_memory[33692] = 3'b111;
        rom_memory[33693] = 3'b111;
        rom_memory[33694] = 3'b111;
        rom_memory[33695] = 3'b111;
        rom_memory[33696] = 3'b111;
        rom_memory[33697] = 3'b111;
        rom_memory[33698] = 3'b111;
        rom_memory[33699] = 3'b110;
        rom_memory[33700] = 3'b110;
        rom_memory[33701] = 3'b110;
        rom_memory[33702] = 3'b110;
        rom_memory[33703] = 3'b110;
        rom_memory[33704] = 3'b110;
        rom_memory[33705] = 3'b110;
        rom_memory[33706] = 3'b110;
        rom_memory[33707] = 3'b110;
        rom_memory[33708] = 3'b110;
        rom_memory[33709] = 3'b110;
        rom_memory[33710] = 3'b110;
        rom_memory[33711] = 3'b110;
        rom_memory[33712] = 3'b110;
        rom_memory[33713] = 3'b110;
        rom_memory[33714] = 3'b110;
        rom_memory[33715] = 3'b110;
        rom_memory[33716] = 3'b110;
        rom_memory[33717] = 3'b110;
        rom_memory[33718] = 3'b110;
        rom_memory[33719] = 3'b110;
        rom_memory[33720] = 3'b110;
        rom_memory[33721] = 3'b110;
        rom_memory[33722] = 3'b110;
        rom_memory[33723] = 3'b110;
        rom_memory[33724] = 3'b110;
        rom_memory[33725] = 3'b110;
        rom_memory[33726] = 3'b110;
        rom_memory[33727] = 3'b110;
        rom_memory[33728] = 3'b110;
        rom_memory[33729] = 3'b110;
        rom_memory[33730] = 3'b110;
        rom_memory[33731] = 3'b110;
        rom_memory[33732] = 3'b110;
        rom_memory[33733] = 3'b110;
        rom_memory[33734] = 3'b110;
        rom_memory[33735] = 3'b110;
        rom_memory[33736] = 3'b110;
        rom_memory[33737] = 3'b110;
        rom_memory[33738] = 3'b110;
        rom_memory[33739] = 3'b000;
        rom_memory[33740] = 3'b000;
        rom_memory[33741] = 3'b000;
        rom_memory[33742] = 3'b000;
        rom_memory[33743] = 3'b000;
        rom_memory[33744] = 3'b000;
        rom_memory[33745] = 3'b111;
        rom_memory[33746] = 3'b100;
        rom_memory[33747] = 3'b000;
        rom_memory[33748] = 3'b100;
        rom_memory[33749] = 3'b110;
        rom_memory[33750] = 3'b000;
        rom_memory[33751] = 3'b000;
        rom_memory[33752] = 3'b000;
        rom_memory[33753] = 3'b100;
        rom_memory[33754] = 3'b110;
        rom_memory[33755] = 3'b110;
        rom_memory[33756] = 3'b110;
        rom_memory[33757] = 3'b110;
        rom_memory[33758] = 3'b110;
        rom_memory[33759] = 3'b110;
        rom_memory[33760] = 3'b110;
        rom_memory[33761] = 3'b110;
        rom_memory[33762] = 3'b110;
        rom_memory[33763] = 3'b110;
        rom_memory[33764] = 3'b110;
        rom_memory[33765] = 3'b110;
        rom_memory[33766] = 3'b110;
        rom_memory[33767] = 3'b110;
        rom_memory[33768] = 3'b110;
        rom_memory[33769] = 3'b110;
        rom_memory[33770] = 3'b110;
        rom_memory[33771] = 3'b110;
        rom_memory[33772] = 3'b110;
        rom_memory[33773] = 3'b110;
        rom_memory[33774] = 3'b110;
        rom_memory[33775] = 3'b110;
        rom_memory[33776] = 3'b110;
        rom_memory[33777] = 3'b110;
        rom_memory[33778] = 3'b110;
        rom_memory[33779] = 3'b110;
        rom_memory[33780] = 3'b110;
        rom_memory[33781] = 3'b110;
        rom_memory[33782] = 3'b110;
        rom_memory[33783] = 3'b110;
        rom_memory[33784] = 3'b110;
        rom_memory[33785] = 3'b110;
        rom_memory[33786] = 3'b111;
        rom_memory[33787] = 3'b110;
        rom_memory[33788] = 3'b111;
        rom_memory[33789] = 3'b111;
        rom_memory[33790] = 3'b111;
        rom_memory[33791] = 3'b111;
        rom_memory[33792] = 3'b111;
        rom_memory[33793] = 3'b111;
        rom_memory[33794] = 3'b111;
        rom_memory[33795] = 3'b111;
        rom_memory[33796] = 3'b111;
        rom_memory[33797] = 3'b111;
        rom_memory[33798] = 3'b111;
        rom_memory[33799] = 3'b111;
        rom_memory[33800] = 3'b111;
        rom_memory[33801] = 3'b111;
        rom_memory[33802] = 3'b111;
        rom_memory[33803] = 3'b111;
        rom_memory[33804] = 3'b111;
        rom_memory[33805] = 3'b111;
        rom_memory[33806] = 3'b111;
        rom_memory[33807] = 3'b111;
        rom_memory[33808] = 3'b111;
        rom_memory[33809] = 3'b111;
        rom_memory[33810] = 3'b111;
        rom_memory[33811] = 3'b111;
        rom_memory[33812] = 3'b111;
        rom_memory[33813] = 3'b111;
        rom_memory[33814] = 3'b111;
        rom_memory[33815] = 3'b111;
        rom_memory[33816] = 3'b111;
        rom_memory[33817] = 3'b111;
        rom_memory[33818] = 3'b111;
        rom_memory[33819] = 3'b111;
        rom_memory[33820] = 3'b111;
        rom_memory[33821] = 3'b111;
        rom_memory[33822] = 3'b111;
        rom_memory[33823] = 3'b111;
        rom_memory[33824] = 3'b111;
        rom_memory[33825] = 3'b111;
        rom_memory[33826] = 3'b111;
        rom_memory[33827] = 3'b111;
        rom_memory[33828] = 3'b111;
        rom_memory[33829] = 3'b111;
        rom_memory[33830] = 3'b111;
        rom_memory[33831] = 3'b111;
        rom_memory[33832] = 3'b111;
        rom_memory[33833] = 3'b111;
        rom_memory[33834] = 3'b111;
        rom_memory[33835] = 3'b111;
        rom_memory[33836] = 3'b111;
        rom_memory[33837] = 3'b111;
        rom_memory[33838] = 3'b111;
        rom_memory[33839] = 3'b111;
        rom_memory[33840] = 3'b110;
        rom_memory[33841] = 3'b110;
        rom_memory[33842] = 3'b110;
        rom_memory[33843] = 3'b110;
        rom_memory[33844] = 3'b110;
        rom_memory[33845] = 3'b111;
        rom_memory[33846] = 3'b111;
        rom_memory[33847] = 3'b111;
        rom_memory[33848] = 3'b111;
        rom_memory[33849] = 3'b111;
        rom_memory[33850] = 3'b111;
        rom_memory[33851] = 3'b111;
        rom_memory[33852] = 3'b111;
        rom_memory[33853] = 3'b111;
        rom_memory[33854] = 3'b111;
        rom_memory[33855] = 3'b111;
        rom_memory[33856] = 3'b111;
        rom_memory[33857] = 3'b111;
        rom_memory[33858] = 3'b111;
        rom_memory[33859] = 3'b111;
        rom_memory[33860] = 3'b111;
        rom_memory[33861] = 3'b110;
        rom_memory[33862] = 3'b110;
        rom_memory[33863] = 3'b110;
        rom_memory[33864] = 3'b111;
        rom_memory[33865] = 3'b111;
        rom_memory[33866] = 3'b111;
        rom_memory[33867] = 3'b111;
        rom_memory[33868] = 3'b111;
        rom_memory[33869] = 3'b111;
        rom_memory[33870] = 3'b111;
        rom_memory[33871] = 3'b111;
        rom_memory[33872] = 3'b111;
        rom_memory[33873] = 3'b111;
        rom_memory[33874] = 3'b110;
        rom_memory[33875] = 3'b110;
        rom_memory[33876] = 3'b110;
        rom_memory[33877] = 3'b110;
        rom_memory[33878] = 3'b110;
        rom_memory[33879] = 3'b110;
        rom_memory[33880] = 3'b110;
        rom_memory[33881] = 3'b110;
        rom_memory[33882] = 3'b110;
        rom_memory[33883] = 3'b110;
        rom_memory[33884] = 3'b110;
        rom_memory[33885] = 3'b110;
        rom_memory[33886] = 3'b111;
        rom_memory[33887] = 3'b111;
        rom_memory[33888] = 3'b111;
        rom_memory[33889] = 3'b111;
        rom_memory[33890] = 3'b111;
        rom_memory[33891] = 3'b111;
        rom_memory[33892] = 3'b111;
        rom_memory[33893] = 3'b111;
        rom_memory[33894] = 3'b111;
        rom_memory[33895] = 3'b111;
        rom_memory[33896] = 3'b111;
        rom_memory[33897] = 3'b111;
        rom_memory[33898] = 3'b111;
        rom_memory[33899] = 3'b111;
        rom_memory[33900] = 3'b111;
        rom_memory[33901] = 3'b111;
        rom_memory[33902] = 3'b000;
        rom_memory[33903] = 3'b000;
        rom_memory[33904] = 3'b000;
        rom_memory[33905] = 3'b000;
        rom_memory[33906] = 3'b000;
        rom_memory[33907] = 3'b000;
        rom_memory[33908] = 3'b000;
        rom_memory[33909] = 3'b000;
        rom_memory[33910] = 3'b000;
        rom_memory[33911] = 3'b000;
        rom_memory[33912] = 3'b000;
        rom_memory[33913] = 3'b111;
        rom_memory[33914] = 3'b100;
        rom_memory[33915] = 3'b000;
        rom_memory[33916] = 3'b000;
        rom_memory[33917] = 3'b111;
        rom_memory[33918] = 3'b000;
        rom_memory[33919] = 3'b000;
        rom_memory[33920] = 3'b000;
        rom_memory[33921] = 3'b000;
        rom_memory[33922] = 3'b000;
        rom_memory[33923] = 3'b000;
        rom_memory[33924] = 3'b000;
        rom_memory[33925] = 3'b000;
        rom_memory[33926] = 3'b000;
        rom_memory[33927] = 3'b000;
        rom_memory[33928] = 3'b100;
        rom_memory[33929] = 3'b100;
        rom_memory[33930] = 3'b110;
        rom_memory[33931] = 3'b111;
        rom_memory[33932] = 3'b111;
        rom_memory[33933] = 3'b110;
        rom_memory[33934] = 3'b111;
        rom_memory[33935] = 3'b111;
        rom_memory[33936] = 3'b111;
        rom_memory[33937] = 3'b111;
        rom_memory[33938] = 3'b111;
        rom_memory[33939] = 3'b110;
        rom_memory[33940] = 3'b110;
        rom_memory[33941] = 3'b110;
        rom_memory[33942] = 3'b110;
        rom_memory[33943] = 3'b110;
        rom_memory[33944] = 3'b110;
        rom_memory[33945] = 3'b110;
        rom_memory[33946] = 3'b110;
        rom_memory[33947] = 3'b110;
        rom_memory[33948] = 3'b110;
        rom_memory[33949] = 3'b110;
        rom_memory[33950] = 3'b110;
        rom_memory[33951] = 3'b110;
        rom_memory[33952] = 3'b110;
        rom_memory[33953] = 3'b110;
        rom_memory[33954] = 3'b110;
        rom_memory[33955] = 3'b110;
        rom_memory[33956] = 3'b110;
        rom_memory[33957] = 3'b110;
        rom_memory[33958] = 3'b110;
        rom_memory[33959] = 3'b110;
        rom_memory[33960] = 3'b110;
        rom_memory[33961] = 3'b110;
        rom_memory[33962] = 3'b110;
        rom_memory[33963] = 3'b110;
        rom_memory[33964] = 3'b110;
        rom_memory[33965] = 3'b110;
        rom_memory[33966] = 3'b110;
        rom_memory[33967] = 3'b110;
        rom_memory[33968] = 3'b110;
        rom_memory[33969] = 3'b110;
        rom_memory[33970] = 3'b110;
        rom_memory[33971] = 3'b110;
        rom_memory[33972] = 3'b110;
        rom_memory[33973] = 3'b110;
        rom_memory[33974] = 3'b110;
        rom_memory[33975] = 3'b110;
        rom_memory[33976] = 3'b110;
        rom_memory[33977] = 3'b110;
        rom_memory[33978] = 3'b110;
        rom_memory[33979] = 3'b111;
        rom_memory[33980] = 3'b000;
        rom_memory[33981] = 3'b000;
        rom_memory[33982] = 3'b000;
        rom_memory[33983] = 3'b000;
        rom_memory[33984] = 3'b000;
        rom_memory[33985] = 3'b000;
        rom_memory[33986] = 3'b111;
        rom_memory[33987] = 3'b100;
        rom_memory[33988] = 3'b000;
        rom_memory[33989] = 3'b100;
        rom_memory[33990] = 3'b110;
        rom_memory[33991] = 3'b000;
        rom_memory[33992] = 3'b000;
        rom_memory[33993] = 3'b000;
        rom_memory[33994] = 3'b100;
        rom_memory[33995] = 3'b111;
        rom_memory[33996] = 3'b110;
        rom_memory[33997] = 3'b110;
        rom_memory[33998] = 3'b110;
        rom_memory[33999] = 3'b110;
        rom_memory[34000] = 3'b110;
        rom_memory[34001] = 3'b110;
        rom_memory[34002] = 3'b110;
        rom_memory[34003] = 3'b110;
        rom_memory[34004] = 3'b110;
        rom_memory[34005] = 3'b110;
        rom_memory[34006] = 3'b110;
        rom_memory[34007] = 3'b110;
        rom_memory[34008] = 3'b110;
        rom_memory[34009] = 3'b110;
        rom_memory[34010] = 3'b110;
        rom_memory[34011] = 3'b110;
        rom_memory[34012] = 3'b110;
        rom_memory[34013] = 3'b110;
        rom_memory[34014] = 3'b110;
        rom_memory[34015] = 3'b110;
        rom_memory[34016] = 3'b110;
        rom_memory[34017] = 3'b110;
        rom_memory[34018] = 3'b110;
        rom_memory[34019] = 3'b110;
        rom_memory[34020] = 3'b110;
        rom_memory[34021] = 3'b110;
        rom_memory[34022] = 3'b110;
        rom_memory[34023] = 3'b110;
        rom_memory[34024] = 3'b110;
        rom_memory[34025] = 3'b110;
        rom_memory[34026] = 3'b110;
        rom_memory[34027] = 3'b110;
        rom_memory[34028] = 3'b111;
        rom_memory[34029] = 3'b111;
        rom_memory[34030] = 3'b111;
        rom_memory[34031] = 3'b111;
        rom_memory[34032] = 3'b111;
        rom_memory[34033] = 3'b111;
        rom_memory[34034] = 3'b111;
        rom_memory[34035] = 3'b111;
        rom_memory[34036] = 3'b111;
        rom_memory[34037] = 3'b111;
        rom_memory[34038] = 3'b111;
        rom_memory[34039] = 3'b111;
        rom_memory[34040] = 3'b111;
        rom_memory[34041] = 3'b111;
        rom_memory[34042] = 3'b111;
        rom_memory[34043] = 3'b111;
        rom_memory[34044] = 3'b111;
        rom_memory[34045] = 3'b111;
        rom_memory[34046] = 3'b111;
        rom_memory[34047] = 3'b111;
        rom_memory[34048] = 3'b111;
        rom_memory[34049] = 3'b111;
        rom_memory[34050] = 3'b111;
        rom_memory[34051] = 3'b111;
        rom_memory[34052] = 3'b111;
        rom_memory[34053] = 3'b111;
        rom_memory[34054] = 3'b111;
        rom_memory[34055] = 3'b111;
        rom_memory[34056] = 3'b111;
        rom_memory[34057] = 3'b111;
        rom_memory[34058] = 3'b111;
        rom_memory[34059] = 3'b111;
        rom_memory[34060] = 3'b111;
        rom_memory[34061] = 3'b111;
        rom_memory[34062] = 3'b111;
        rom_memory[34063] = 3'b111;
        rom_memory[34064] = 3'b111;
        rom_memory[34065] = 3'b111;
        rom_memory[34066] = 3'b111;
        rom_memory[34067] = 3'b111;
        rom_memory[34068] = 3'b111;
        rom_memory[34069] = 3'b111;
        rom_memory[34070] = 3'b111;
        rom_memory[34071] = 3'b111;
        rom_memory[34072] = 3'b111;
        rom_memory[34073] = 3'b111;
        rom_memory[34074] = 3'b111;
        rom_memory[34075] = 3'b111;
        rom_memory[34076] = 3'b111;
        rom_memory[34077] = 3'b111;
        rom_memory[34078] = 3'b111;
        rom_memory[34079] = 3'b111;
        rom_memory[34080] = 3'b110;
        rom_memory[34081] = 3'b110;
        rom_memory[34082] = 3'b110;
        rom_memory[34083] = 3'b110;
        rom_memory[34084] = 3'b110;
        rom_memory[34085] = 3'b111;
        rom_memory[34086] = 3'b111;
        rom_memory[34087] = 3'b111;
        rom_memory[34088] = 3'b111;
        rom_memory[34089] = 3'b111;
        rom_memory[34090] = 3'b111;
        rom_memory[34091] = 3'b111;
        rom_memory[34092] = 3'b111;
        rom_memory[34093] = 3'b111;
        rom_memory[34094] = 3'b111;
        rom_memory[34095] = 3'b111;
        rom_memory[34096] = 3'b111;
        rom_memory[34097] = 3'b111;
        rom_memory[34098] = 3'b111;
        rom_memory[34099] = 3'b111;
        rom_memory[34100] = 3'b111;
        rom_memory[34101] = 3'b111;
        rom_memory[34102] = 3'b110;
        rom_memory[34103] = 3'b110;
        rom_memory[34104] = 3'b111;
        rom_memory[34105] = 3'b111;
        rom_memory[34106] = 3'b111;
        rom_memory[34107] = 3'b111;
        rom_memory[34108] = 3'b111;
        rom_memory[34109] = 3'b111;
        rom_memory[34110] = 3'b111;
        rom_memory[34111] = 3'b111;
        rom_memory[34112] = 3'b111;
        rom_memory[34113] = 3'b110;
        rom_memory[34114] = 3'b110;
        rom_memory[34115] = 3'b110;
        rom_memory[34116] = 3'b110;
        rom_memory[34117] = 3'b110;
        rom_memory[34118] = 3'b110;
        rom_memory[34119] = 3'b110;
        rom_memory[34120] = 3'b110;
        rom_memory[34121] = 3'b110;
        rom_memory[34122] = 3'b110;
        rom_memory[34123] = 3'b110;
        rom_memory[34124] = 3'b110;
        rom_memory[34125] = 3'b110;
        rom_memory[34126] = 3'b111;
        rom_memory[34127] = 3'b111;
        rom_memory[34128] = 3'b111;
        rom_memory[34129] = 3'b111;
        rom_memory[34130] = 3'b111;
        rom_memory[34131] = 3'b111;
        rom_memory[34132] = 3'b111;
        rom_memory[34133] = 3'b111;
        rom_memory[34134] = 3'b111;
        rom_memory[34135] = 3'b111;
        rom_memory[34136] = 3'b111;
        rom_memory[34137] = 3'b111;
        rom_memory[34138] = 3'b111;
        rom_memory[34139] = 3'b111;
        rom_memory[34140] = 3'b111;
        rom_memory[34141] = 3'b111;
        rom_memory[34142] = 3'b111;
        rom_memory[34143] = 3'b000;
        rom_memory[34144] = 3'b000;
        rom_memory[34145] = 3'b000;
        rom_memory[34146] = 3'b000;
        rom_memory[34147] = 3'b000;
        rom_memory[34148] = 3'b000;
        rom_memory[34149] = 3'b000;
        rom_memory[34150] = 3'b000;
        rom_memory[34151] = 3'b000;
        rom_memory[34152] = 3'b111;
        rom_memory[34153] = 3'b000;
        rom_memory[34154] = 3'b000;
        rom_memory[34155] = 3'b000;
        rom_memory[34156] = 3'b100;
        rom_memory[34157] = 3'b110;
        rom_memory[34158] = 3'b000;
        rom_memory[34159] = 3'b000;
        rom_memory[34160] = 3'b000;
        rom_memory[34161] = 3'b110;
        rom_memory[34162] = 3'b000;
        rom_memory[34163] = 3'b000;
        rom_memory[34164] = 3'b000;
        rom_memory[34165] = 3'b000;
        rom_memory[34166] = 3'b000;
        rom_memory[34167] = 3'b000;
        rom_memory[34168] = 3'b000;
        rom_memory[34169] = 3'b100;
        rom_memory[34170] = 3'b100;
        rom_memory[34171] = 3'b111;
        rom_memory[34172] = 3'b111;
        rom_memory[34173] = 3'b110;
        rom_memory[34174] = 3'b110;
        rom_memory[34175] = 3'b111;
        rom_memory[34176] = 3'b111;
        rom_memory[34177] = 3'b111;
        rom_memory[34178] = 3'b110;
        rom_memory[34179] = 3'b110;
        rom_memory[34180] = 3'b110;
        rom_memory[34181] = 3'b110;
        rom_memory[34182] = 3'b110;
        rom_memory[34183] = 3'b110;
        rom_memory[34184] = 3'b110;
        rom_memory[34185] = 3'b110;
        rom_memory[34186] = 3'b110;
        rom_memory[34187] = 3'b110;
        rom_memory[34188] = 3'b110;
        rom_memory[34189] = 3'b110;
        rom_memory[34190] = 3'b110;
        rom_memory[34191] = 3'b110;
        rom_memory[34192] = 3'b110;
        rom_memory[34193] = 3'b110;
        rom_memory[34194] = 3'b110;
        rom_memory[34195] = 3'b110;
        rom_memory[34196] = 3'b110;
        rom_memory[34197] = 3'b110;
        rom_memory[34198] = 3'b110;
        rom_memory[34199] = 3'b110;
        rom_memory[34200] = 3'b110;
        rom_memory[34201] = 3'b110;
        rom_memory[34202] = 3'b110;
        rom_memory[34203] = 3'b110;
        rom_memory[34204] = 3'b110;
        rom_memory[34205] = 3'b110;
        rom_memory[34206] = 3'b110;
        rom_memory[34207] = 3'b110;
        rom_memory[34208] = 3'b110;
        rom_memory[34209] = 3'b110;
        rom_memory[34210] = 3'b110;
        rom_memory[34211] = 3'b110;
        rom_memory[34212] = 3'b110;
        rom_memory[34213] = 3'b110;
        rom_memory[34214] = 3'b110;
        rom_memory[34215] = 3'b110;
        rom_memory[34216] = 3'b110;
        rom_memory[34217] = 3'b110;
        rom_memory[34218] = 3'b110;
        rom_memory[34219] = 3'b110;
        rom_memory[34220] = 3'b110;
        rom_memory[34221] = 3'b100;
        rom_memory[34222] = 3'b000;
        rom_memory[34223] = 3'b000;
        rom_memory[34224] = 3'b000;
        rom_memory[34225] = 3'b000;
        rom_memory[34226] = 3'b000;
        rom_memory[34227] = 3'b111;
        rom_memory[34228] = 3'b110;
        rom_memory[34229] = 3'b000;
        rom_memory[34230] = 3'b100;
        rom_memory[34231] = 3'b110;
        rom_memory[34232] = 3'b100;
        rom_memory[34233] = 3'b000;
        rom_memory[34234] = 3'b000;
        rom_memory[34235] = 3'b100;
        rom_memory[34236] = 3'b110;
        rom_memory[34237] = 3'b110;
        rom_memory[34238] = 3'b110;
        rom_memory[34239] = 3'b110;
        rom_memory[34240] = 3'b110;
        rom_memory[34241] = 3'b110;
        rom_memory[34242] = 3'b110;
        rom_memory[34243] = 3'b110;
        rom_memory[34244] = 3'b110;
        rom_memory[34245] = 3'b110;
        rom_memory[34246] = 3'b110;
        rom_memory[34247] = 3'b110;
        rom_memory[34248] = 3'b110;
        rom_memory[34249] = 3'b110;
        rom_memory[34250] = 3'b110;
        rom_memory[34251] = 3'b110;
        rom_memory[34252] = 3'b110;
        rom_memory[34253] = 3'b110;
        rom_memory[34254] = 3'b110;
        rom_memory[34255] = 3'b110;
        rom_memory[34256] = 3'b110;
        rom_memory[34257] = 3'b110;
        rom_memory[34258] = 3'b110;
        rom_memory[34259] = 3'b110;
        rom_memory[34260] = 3'b110;
        rom_memory[34261] = 3'b110;
        rom_memory[34262] = 3'b110;
        rom_memory[34263] = 3'b110;
        rom_memory[34264] = 3'b110;
        rom_memory[34265] = 3'b110;
        rom_memory[34266] = 3'b110;
        rom_memory[34267] = 3'b110;
        rom_memory[34268] = 3'b110;
        rom_memory[34269] = 3'b111;
        rom_memory[34270] = 3'b111;
        rom_memory[34271] = 3'b111;
        rom_memory[34272] = 3'b111;
        rom_memory[34273] = 3'b111;
        rom_memory[34274] = 3'b111;
        rom_memory[34275] = 3'b111;
        rom_memory[34276] = 3'b111;
        rom_memory[34277] = 3'b111;
        rom_memory[34278] = 3'b111;
        rom_memory[34279] = 3'b111;
        rom_memory[34280] = 3'b111;
        rom_memory[34281] = 3'b111;
        rom_memory[34282] = 3'b111;
        rom_memory[34283] = 3'b111;
        rom_memory[34284] = 3'b111;
        rom_memory[34285] = 3'b111;
        rom_memory[34286] = 3'b111;
        rom_memory[34287] = 3'b111;
        rom_memory[34288] = 3'b111;
        rom_memory[34289] = 3'b111;
        rom_memory[34290] = 3'b111;
        rom_memory[34291] = 3'b111;
        rom_memory[34292] = 3'b111;
        rom_memory[34293] = 3'b111;
        rom_memory[34294] = 3'b111;
        rom_memory[34295] = 3'b111;
        rom_memory[34296] = 3'b111;
        rom_memory[34297] = 3'b111;
        rom_memory[34298] = 3'b111;
        rom_memory[34299] = 3'b111;
        rom_memory[34300] = 3'b111;
        rom_memory[34301] = 3'b111;
        rom_memory[34302] = 3'b111;
        rom_memory[34303] = 3'b111;
        rom_memory[34304] = 3'b111;
        rom_memory[34305] = 3'b111;
        rom_memory[34306] = 3'b111;
        rom_memory[34307] = 3'b111;
        rom_memory[34308] = 3'b111;
        rom_memory[34309] = 3'b111;
        rom_memory[34310] = 3'b111;
        rom_memory[34311] = 3'b111;
        rom_memory[34312] = 3'b111;
        rom_memory[34313] = 3'b111;
        rom_memory[34314] = 3'b111;
        rom_memory[34315] = 3'b111;
        rom_memory[34316] = 3'b111;
        rom_memory[34317] = 3'b111;
        rom_memory[34318] = 3'b111;
        rom_memory[34319] = 3'b111;
        rom_memory[34320] = 3'b110;
        rom_memory[34321] = 3'b110;
        rom_memory[34322] = 3'b110;
        rom_memory[34323] = 3'b110;
        rom_memory[34324] = 3'b110;
        rom_memory[34325] = 3'b111;
        rom_memory[34326] = 3'b111;
        rom_memory[34327] = 3'b111;
        rom_memory[34328] = 3'b111;
        rom_memory[34329] = 3'b111;
        rom_memory[34330] = 3'b111;
        rom_memory[34331] = 3'b111;
        rom_memory[34332] = 3'b111;
        rom_memory[34333] = 3'b111;
        rom_memory[34334] = 3'b111;
        rom_memory[34335] = 3'b111;
        rom_memory[34336] = 3'b111;
        rom_memory[34337] = 3'b111;
        rom_memory[34338] = 3'b111;
        rom_memory[34339] = 3'b111;
        rom_memory[34340] = 3'b111;
        rom_memory[34341] = 3'b111;
        rom_memory[34342] = 3'b110;
        rom_memory[34343] = 3'b110;
        rom_memory[34344] = 3'b110;
        rom_memory[34345] = 3'b111;
        rom_memory[34346] = 3'b111;
        rom_memory[34347] = 3'b111;
        rom_memory[34348] = 3'b111;
        rom_memory[34349] = 3'b111;
        rom_memory[34350] = 3'b111;
        rom_memory[34351] = 3'b111;
        rom_memory[34352] = 3'b111;
        rom_memory[34353] = 3'b110;
        rom_memory[34354] = 3'b110;
        rom_memory[34355] = 3'b110;
        rom_memory[34356] = 3'b110;
        rom_memory[34357] = 3'b110;
        rom_memory[34358] = 3'b110;
        rom_memory[34359] = 3'b110;
        rom_memory[34360] = 3'b110;
        rom_memory[34361] = 3'b110;
        rom_memory[34362] = 3'b110;
        rom_memory[34363] = 3'b110;
        rom_memory[34364] = 3'b110;
        rom_memory[34365] = 3'b110;
        rom_memory[34366] = 3'b111;
        rom_memory[34367] = 3'b111;
        rom_memory[34368] = 3'b111;
        rom_memory[34369] = 3'b111;
        rom_memory[34370] = 3'b111;
        rom_memory[34371] = 3'b111;
        rom_memory[34372] = 3'b111;
        rom_memory[34373] = 3'b111;
        rom_memory[34374] = 3'b111;
        rom_memory[34375] = 3'b111;
        rom_memory[34376] = 3'b111;
        rom_memory[34377] = 3'b111;
        rom_memory[34378] = 3'b111;
        rom_memory[34379] = 3'b111;
        rom_memory[34380] = 3'b111;
        rom_memory[34381] = 3'b111;
        rom_memory[34382] = 3'b111;
        rom_memory[34383] = 3'b000;
        rom_memory[34384] = 3'b000;
        rom_memory[34385] = 3'b000;
        rom_memory[34386] = 3'b000;
        rom_memory[34387] = 3'b000;
        rom_memory[34388] = 3'b000;
        rom_memory[34389] = 3'b000;
        rom_memory[34390] = 3'b000;
        rom_memory[34391] = 3'b000;
        rom_memory[34392] = 3'b000;
        rom_memory[34393] = 3'b000;
        rom_memory[34394] = 3'b000;
        rom_memory[34395] = 3'b000;
        rom_memory[34396] = 3'b000;
        rom_memory[34397] = 3'b100;
        rom_memory[34398] = 3'b000;
        rom_memory[34399] = 3'b000;
        rom_memory[34400] = 3'b100;
        rom_memory[34401] = 3'b110;
        rom_memory[34402] = 3'b000;
        rom_memory[34403] = 3'b000;
        rom_memory[34404] = 3'b000;
        rom_memory[34405] = 3'b000;
        rom_memory[34406] = 3'b000;
        rom_memory[34407] = 3'b000;
        rom_memory[34408] = 3'b000;
        rom_memory[34409] = 3'b100;
        rom_memory[34410] = 3'b000;
        rom_memory[34411] = 3'b111;
        rom_memory[34412] = 3'b111;
        rom_memory[34413] = 3'b110;
        rom_memory[34414] = 3'b110;
        rom_memory[34415] = 3'b111;
        rom_memory[34416] = 3'b111;
        rom_memory[34417] = 3'b111;
        rom_memory[34418] = 3'b110;
        rom_memory[34419] = 3'b110;
        rom_memory[34420] = 3'b110;
        rom_memory[34421] = 3'b110;
        rom_memory[34422] = 3'b110;
        rom_memory[34423] = 3'b110;
        rom_memory[34424] = 3'b110;
        rom_memory[34425] = 3'b110;
        rom_memory[34426] = 3'b110;
        rom_memory[34427] = 3'b110;
        rom_memory[34428] = 3'b110;
        rom_memory[34429] = 3'b110;
        rom_memory[34430] = 3'b110;
        rom_memory[34431] = 3'b110;
        rom_memory[34432] = 3'b110;
        rom_memory[34433] = 3'b110;
        rom_memory[34434] = 3'b110;
        rom_memory[34435] = 3'b110;
        rom_memory[34436] = 3'b110;
        rom_memory[34437] = 3'b110;
        rom_memory[34438] = 3'b110;
        rom_memory[34439] = 3'b110;
        rom_memory[34440] = 3'b110;
        rom_memory[34441] = 3'b110;
        rom_memory[34442] = 3'b110;
        rom_memory[34443] = 3'b110;
        rom_memory[34444] = 3'b110;
        rom_memory[34445] = 3'b110;
        rom_memory[34446] = 3'b110;
        rom_memory[34447] = 3'b110;
        rom_memory[34448] = 3'b110;
        rom_memory[34449] = 3'b110;
        rom_memory[34450] = 3'b110;
        rom_memory[34451] = 3'b110;
        rom_memory[34452] = 3'b110;
        rom_memory[34453] = 3'b110;
        rom_memory[34454] = 3'b110;
        rom_memory[34455] = 3'b110;
        rom_memory[34456] = 3'b110;
        rom_memory[34457] = 3'b110;
        rom_memory[34458] = 3'b110;
        rom_memory[34459] = 3'b110;
        rom_memory[34460] = 3'b110;
        rom_memory[34461] = 3'b110;
        rom_memory[34462] = 3'b110;
        rom_memory[34463] = 3'b000;
        rom_memory[34464] = 3'b000;
        rom_memory[34465] = 3'b000;
        rom_memory[34466] = 3'b000;
        rom_memory[34467] = 3'b000;
        rom_memory[34468] = 3'b111;
        rom_memory[34469] = 3'b110;
        rom_memory[34470] = 3'b000;
        rom_memory[34471] = 3'b100;
        rom_memory[34472] = 3'b110;
        rom_memory[34473] = 3'b100;
        rom_memory[34474] = 3'b000;
        rom_memory[34475] = 3'b000;
        rom_memory[34476] = 3'b100;
        rom_memory[34477] = 3'b110;
        rom_memory[34478] = 3'b110;
        rom_memory[34479] = 3'b110;
        rom_memory[34480] = 3'b110;
        rom_memory[34481] = 3'b110;
        rom_memory[34482] = 3'b110;
        rom_memory[34483] = 3'b110;
        rom_memory[34484] = 3'b110;
        rom_memory[34485] = 3'b110;
        rom_memory[34486] = 3'b110;
        rom_memory[34487] = 3'b110;
        rom_memory[34488] = 3'b110;
        rom_memory[34489] = 3'b110;
        rom_memory[34490] = 3'b110;
        rom_memory[34491] = 3'b110;
        rom_memory[34492] = 3'b110;
        rom_memory[34493] = 3'b110;
        rom_memory[34494] = 3'b110;
        rom_memory[34495] = 3'b110;
        rom_memory[34496] = 3'b110;
        rom_memory[34497] = 3'b110;
        rom_memory[34498] = 3'b110;
        rom_memory[34499] = 3'b110;
        rom_memory[34500] = 3'b110;
        rom_memory[34501] = 3'b110;
        rom_memory[34502] = 3'b110;
        rom_memory[34503] = 3'b110;
        rom_memory[34504] = 3'b110;
        rom_memory[34505] = 3'b110;
        rom_memory[34506] = 3'b110;
        rom_memory[34507] = 3'b110;
        rom_memory[34508] = 3'b110;
        rom_memory[34509] = 3'b111;
        rom_memory[34510] = 3'b111;
        rom_memory[34511] = 3'b111;
        rom_memory[34512] = 3'b111;
        rom_memory[34513] = 3'b111;
        rom_memory[34514] = 3'b111;
        rom_memory[34515] = 3'b111;
        rom_memory[34516] = 3'b111;
        rom_memory[34517] = 3'b111;
        rom_memory[34518] = 3'b111;
        rom_memory[34519] = 3'b111;
        rom_memory[34520] = 3'b111;
        rom_memory[34521] = 3'b111;
        rom_memory[34522] = 3'b111;
        rom_memory[34523] = 3'b111;
        rom_memory[34524] = 3'b111;
        rom_memory[34525] = 3'b111;
        rom_memory[34526] = 3'b111;
        rom_memory[34527] = 3'b111;
        rom_memory[34528] = 3'b111;
        rom_memory[34529] = 3'b111;
        rom_memory[34530] = 3'b111;
        rom_memory[34531] = 3'b111;
        rom_memory[34532] = 3'b111;
        rom_memory[34533] = 3'b111;
        rom_memory[34534] = 3'b111;
        rom_memory[34535] = 3'b111;
        rom_memory[34536] = 3'b111;
        rom_memory[34537] = 3'b111;
        rom_memory[34538] = 3'b111;
        rom_memory[34539] = 3'b111;
        rom_memory[34540] = 3'b111;
        rom_memory[34541] = 3'b111;
        rom_memory[34542] = 3'b111;
        rom_memory[34543] = 3'b111;
        rom_memory[34544] = 3'b111;
        rom_memory[34545] = 3'b111;
        rom_memory[34546] = 3'b111;
        rom_memory[34547] = 3'b111;
        rom_memory[34548] = 3'b111;
        rom_memory[34549] = 3'b111;
        rom_memory[34550] = 3'b111;
        rom_memory[34551] = 3'b111;
        rom_memory[34552] = 3'b111;
        rom_memory[34553] = 3'b111;
        rom_memory[34554] = 3'b111;
        rom_memory[34555] = 3'b111;
        rom_memory[34556] = 3'b111;
        rom_memory[34557] = 3'b111;
        rom_memory[34558] = 3'b111;
        rom_memory[34559] = 3'b111;
        rom_memory[34560] = 3'b110;
        rom_memory[34561] = 3'b110;
        rom_memory[34562] = 3'b110;
        rom_memory[34563] = 3'b110;
        rom_memory[34564] = 3'b110;
        rom_memory[34565] = 3'b111;
        rom_memory[34566] = 3'b111;
        rom_memory[34567] = 3'b111;
        rom_memory[34568] = 3'b111;
        rom_memory[34569] = 3'b111;
        rom_memory[34570] = 3'b111;
        rom_memory[34571] = 3'b111;
        rom_memory[34572] = 3'b111;
        rom_memory[34573] = 3'b111;
        rom_memory[34574] = 3'b111;
        rom_memory[34575] = 3'b111;
        rom_memory[34576] = 3'b111;
        rom_memory[34577] = 3'b111;
        rom_memory[34578] = 3'b111;
        rom_memory[34579] = 3'b111;
        rom_memory[34580] = 3'b111;
        rom_memory[34581] = 3'b111;
        rom_memory[34582] = 3'b111;
        rom_memory[34583] = 3'b110;
        rom_memory[34584] = 3'b110;
        rom_memory[34585] = 3'b110;
        rom_memory[34586] = 3'b111;
        rom_memory[34587] = 3'b111;
        rom_memory[34588] = 3'b111;
        rom_memory[34589] = 3'b111;
        rom_memory[34590] = 3'b111;
        rom_memory[34591] = 3'b111;
        rom_memory[34592] = 3'b111;
        rom_memory[34593] = 3'b110;
        rom_memory[34594] = 3'b110;
        rom_memory[34595] = 3'b110;
        rom_memory[34596] = 3'b110;
        rom_memory[34597] = 3'b110;
        rom_memory[34598] = 3'b110;
        rom_memory[34599] = 3'b110;
        rom_memory[34600] = 3'b110;
        rom_memory[34601] = 3'b110;
        rom_memory[34602] = 3'b110;
        rom_memory[34603] = 3'b110;
        rom_memory[34604] = 3'b110;
        rom_memory[34605] = 3'b110;
        rom_memory[34606] = 3'b111;
        rom_memory[34607] = 3'b111;
        rom_memory[34608] = 3'b111;
        rom_memory[34609] = 3'b111;
        rom_memory[34610] = 3'b111;
        rom_memory[34611] = 3'b111;
        rom_memory[34612] = 3'b111;
        rom_memory[34613] = 3'b111;
        rom_memory[34614] = 3'b111;
        rom_memory[34615] = 3'b111;
        rom_memory[34616] = 3'b111;
        rom_memory[34617] = 3'b111;
        rom_memory[34618] = 3'b111;
        rom_memory[34619] = 3'b111;
        rom_memory[34620] = 3'b111;
        rom_memory[34621] = 3'b111;
        rom_memory[34622] = 3'b111;
        rom_memory[34623] = 3'b000;
        rom_memory[34624] = 3'b000;
        rom_memory[34625] = 3'b000;
        rom_memory[34626] = 3'b000;
        rom_memory[34627] = 3'b000;
        rom_memory[34628] = 3'b000;
        rom_memory[34629] = 3'b000;
        rom_memory[34630] = 3'b000;
        rom_memory[34631] = 3'b001;
        rom_memory[34632] = 3'b000;
        rom_memory[34633] = 3'b000;
        rom_memory[34634] = 3'b000;
        rom_memory[34635] = 3'b000;
        rom_memory[34636] = 3'b000;
        rom_memory[34637] = 3'b000;
        rom_memory[34638] = 3'b000;
        rom_memory[34639] = 3'b000;
        rom_memory[34640] = 3'b100;
        rom_memory[34641] = 3'b100;
        rom_memory[34642] = 3'b100;
        rom_memory[34643] = 3'b000;
        rom_memory[34644] = 3'b000;
        rom_memory[34645] = 3'b000;
        rom_memory[34646] = 3'b000;
        rom_memory[34647] = 3'b000;
        rom_memory[34648] = 3'b100;
        rom_memory[34649] = 3'b110;
        rom_memory[34650] = 3'b000;
        rom_memory[34651] = 3'b111;
        rom_memory[34652] = 3'b110;
        rom_memory[34653] = 3'b110;
        rom_memory[34654] = 3'b110;
        rom_memory[34655] = 3'b111;
        rom_memory[34656] = 3'b111;
        rom_memory[34657] = 3'b111;
        rom_memory[34658] = 3'b110;
        rom_memory[34659] = 3'b110;
        rom_memory[34660] = 3'b110;
        rom_memory[34661] = 3'b110;
        rom_memory[34662] = 3'b110;
        rom_memory[34663] = 3'b110;
        rom_memory[34664] = 3'b110;
        rom_memory[34665] = 3'b110;
        rom_memory[34666] = 3'b110;
        rom_memory[34667] = 3'b110;
        rom_memory[34668] = 3'b110;
        rom_memory[34669] = 3'b110;
        rom_memory[34670] = 3'b110;
        rom_memory[34671] = 3'b110;
        rom_memory[34672] = 3'b110;
        rom_memory[34673] = 3'b110;
        rom_memory[34674] = 3'b110;
        rom_memory[34675] = 3'b110;
        rom_memory[34676] = 3'b110;
        rom_memory[34677] = 3'b110;
        rom_memory[34678] = 3'b110;
        rom_memory[34679] = 3'b110;
        rom_memory[34680] = 3'b110;
        rom_memory[34681] = 3'b110;
        rom_memory[34682] = 3'b110;
        rom_memory[34683] = 3'b110;
        rom_memory[34684] = 3'b110;
        rom_memory[34685] = 3'b110;
        rom_memory[34686] = 3'b110;
        rom_memory[34687] = 3'b110;
        rom_memory[34688] = 3'b110;
        rom_memory[34689] = 3'b110;
        rom_memory[34690] = 3'b110;
        rom_memory[34691] = 3'b110;
        rom_memory[34692] = 3'b110;
        rom_memory[34693] = 3'b110;
        rom_memory[34694] = 3'b110;
        rom_memory[34695] = 3'b110;
        rom_memory[34696] = 3'b110;
        rom_memory[34697] = 3'b110;
        rom_memory[34698] = 3'b110;
        rom_memory[34699] = 3'b110;
        rom_memory[34700] = 3'b110;
        rom_memory[34701] = 3'b110;
        rom_memory[34702] = 3'b110;
        rom_memory[34703] = 3'b110;
        rom_memory[34704] = 3'b000;
        rom_memory[34705] = 3'b000;
        rom_memory[34706] = 3'b000;
        rom_memory[34707] = 3'b000;
        rom_memory[34708] = 3'b000;
        rom_memory[34709] = 3'b111;
        rom_memory[34710] = 3'b110;
        rom_memory[34711] = 3'b000;
        rom_memory[34712] = 3'b100;
        rom_memory[34713] = 3'b110;
        rom_memory[34714] = 3'b100;
        rom_memory[34715] = 3'b000;
        rom_memory[34716] = 3'b000;
        rom_memory[34717] = 3'b100;
        rom_memory[34718] = 3'b110;
        rom_memory[34719] = 3'b111;
        rom_memory[34720] = 3'b110;
        rom_memory[34721] = 3'b110;
        rom_memory[34722] = 3'b110;
        rom_memory[34723] = 3'b110;
        rom_memory[34724] = 3'b110;
        rom_memory[34725] = 3'b110;
        rom_memory[34726] = 3'b110;
        rom_memory[34727] = 3'b110;
        rom_memory[34728] = 3'b110;
        rom_memory[34729] = 3'b110;
        rom_memory[34730] = 3'b110;
        rom_memory[34731] = 3'b110;
        rom_memory[34732] = 3'b110;
        rom_memory[34733] = 3'b110;
        rom_memory[34734] = 3'b110;
        rom_memory[34735] = 3'b110;
        rom_memory[34736] = 3'b110;
        rom_memory[34737] = 3'b110;
        rom_memory[34738] = 3'b110;
        rom_memory[34739] = 3'b110;
        rom_memory[34740] = 3'b110;
        rom_memory[34741] = 3'b110;
        rom_memory[34742] = 3'b110;
        rom_memory[34743] = 3'b110;
        rom_memory[34744] = 3'b110;
        rom_memory[34745] = 3'b110;
        rom_memory[34746] = 3'b110;
        rom_memory[34747] = 3'b110;
        rom_memory[34748] = 3'b110;
        rom_memory[34749] = 3'b110;
        rom_memory[34750] = 3'b110;
        rom_memory[34751] = 3'b111;
        rom_memory[34752] = 3'b111;
        rom_memory[34753] = 3'b111;
        rom_memory[34754] = 3'b111;
        rom_memory[34755] = 3'b111;
        rom_memory[34756] = 3'b111;
        rom_memory[34757] = 3'b111;
        rom_memory[34758] = 3'b111;
        rom_memory[34759] = 3'b111;
        rom_memory[34760] = 3'b111;
        rom_memory[34761] = 3'b111;
        rom_memory[34762] = 3'b111;
        rom_memory[34763] = 3'b111;
        rom_memory[34764] = 3'b111;
        rom_memory[34765] = 3'b111;
        rom_memory[34766] = 3'b111;
        rom_memory[34767] = 3'b111;
        rom_memory[34768] = 3'b111;
        rom_memory[34769] = 3'b111;
        rom_memory[34770] = 3'b111;
        rom_memory[34771] = 3'b111;
        rom_memory[34772] = 3'b111;
        rom_memory[34773] = 3'b111;
        rom_memory[34774] = 3'b111;
        rom_memory[34775] = 3'b111;
        rom_memory[34776] = 3'b111;
        rom_memory[34777] = 3'b111;
        rom_memory[34778] = 3'b111;
        rom_memory[34779] = 3'b111;
        rom_memory[34780] = 3'b111;
        rom_memory[34781] = 3'b111;
        rom_memory[34782] = 3'b111;
        rom_memory[34783] = 3'b111;
        rom_memory[34784] = 3'b111;
        rom_memory[34785] = 3'b111;
        rom_memory[34786] = 3'b111;
        rom_memory[34787] = 3'b111;
        rom_memory[34788] = 3'b111;
        rom_memory[34789] = 3'b111;
        rom_memory[34790] = 3'b111;
        rom_memory[34791] = 3'b111;
        rom_memory[34792] = 3'b111;
        rom_memory[34793] = 3'b111;
        rom_memory[34794] = 3'b111;
        rom_memory[34795] = 3'b111;
        rom_memory[34796] = 3'b111;
        rom_memory[34797] = 3'b111;
        rom_memory[34798] = 3'b111;
        rom_memory[34799] = 3'b111;
        rom_memory[34800] = 3'b110;
        rom_memory[34801] = 3'b110;
        rom_memory[34802] = 3'b110;
        rom_memory[34803] = 3'b110;
        rom_memory[34804] = 3'b110;
        rom_memory[34805] = 3'b111;
        rom_memory[34806] = 3'b111;
        rom_memory[34807] = 3'b111;
        rom_memory[34808] = 3'b111;
        rom_memory[34809] = 3'b111;
        rom_memory[34810] = 3'b111;
        rom_memory[34811] = 3'b111;
        rom_memory[34812] = 3'b111;
        rom_memory[34813] = 3'b111;
        rom_memory[34814] = 3'b111;
        rom_memory[34815] = 3'b111;
        rom_memory[34816] = 3'b111;
        rom_memory[34817] = 3'b111;
        rom_memory[34818] = 3'b111;
        rom_memory[34819] = 3'b111;
        rom_memory[34820] = 3'b111;
        rom_memory[34821] = 3'b111;
        rom_memory[34822] = 3'b110;
        rom_memory[34823] = 3'b110;
        rom_memory[34824] = 3'b110;
        rom_memory[34825] = 3'b110;
        rom_memory[34826] = 3'b110;
        rom_memory[34827] = 3'b111;
        rom_memory[34828] = 3'b111;
        rom_memory[34829] = 3'b111;
        rom_memory[34830] = 3'b111;
        rom_memory[34831] = 3'b111;
        rom_memory[34832] = 3'b110;
        rom_memory[34833] = 3'b110;
        rom_memory[34834] = 3'b110;
        rom_memory[34835] = 3'b110;
        rom_memory[34836] = 3'b110;
        rom_memory[34837] = 3'b110;
        rom_memory[34838] = 3'b110;
        rom_memory[34839] = 3'b110;
        rom_memory[34840] = 3'b110;
        rom_memory[34841] = 3'b110;
        rom_memory[34842] = 3'b110;
        rom_memory[34843] = 3'b110;
        rom_memory[34844] = 3'b110;
        rom_memory[34845] = 3'b111;
        rom_memory[34846] = 3'b111;
        rom_memory[34847] = 3'b111;
        rom_memory[34848] = 3'b111;
        rom_memory[34849] = 3'b111;
        rom_memory[34850] = 3'b111;
        rom_memory[34851] = 3'b111;
        rom_memory[34852] = 3'b111;
        rom_memory[34853] = 3'b111;
        rom_memory[34854] = 3'b111;
        rom_memory[34855] = 3'b111;
        rom_memory[34856] = 3'b111;
        rom_memory[34857] = 3'b111;
        rom_memory[34858] = 3'b111;
        rom_memory[34859] = 3'b111;
        rom_memory[34860] = 3'b111;
        rom_memory[34861] = 3'b111;
        rom_memory[34862] = 3'b111;
        rom_memory[34863] = 3'b000;
        rom_memory[34864] = 3'b000;
        rom_memory[34865] = 3'b000;
        rom_memory[34866] = 3'b000;
        rom_memory[34867] = 3'b000;
        rom_memory[34868] = 3'b111;
        rom_memory[34869] = 3'b000;
        rom_memory[34870] = 3'b000;
        rom_memory[34871] = 3'b000;
        rom_memory[34872] = 3'b000;
        rom_memory[34873] = 3'b000;
        rom_memory[34874] = 3'b000;
        rom_memory[34875] = 3'b000;
        rom_memory[34876] = 3'b000;
        rom_memory[34877] = 3'b000;
        rom_memory[34878] = 3'b000;
        rom_memory[34879] = 3'b100;
        rom_memory[34880] = 3'b110;
        rom_memory[34881] = 3'b100;
        rom_memory[34882] = 3'b111;
        rom_memory[34883] = 3'b000;
        rom_memory[34884] = 3'b000;
        rom_memory[34885] = 3'b000;
        rom_memory[34886] = 3'b000;
        rom_memory[34887] = 3'b100;
        rom_memory[34888] = 3'b110;
        rom_memory[34889] = 3'b111;
        rom_memory[34890] = 3'b111;
        rom_memory[34891] = 3'b111;
        rom_memory[34892] = 3'b110;
        rom_memory[34893] = 3'b111;
        rom_memory[34894] = 3'b111;
        rom_memory[34895] = 3'b110;
        rom_memory[34896] = 3'b111;
        rom_memory[34897] = 3'b111;
        rom_memory[34898] = 3'b111;
        rom_memory[34899] = 3'b110;
        rom_memory[34900] = 3'b110;
        rom_memory[34901] = 3'b110;
        rom_memory[34902] = 3'b110;
        rom_memory[34903] = 3'b110;
        rom_memory[34904] = 3'b110;
        rom_memory[34905] = 3'b110;
        rom_memory[34906] = 3'b110;
        rom_memory[34907] = 3'b110;
        rom_memory[34908] = 3'b110;
        rom_memory[34909] = 3'b110;
        rom_memory[34910] = 3'b110;
        rom_memory[34911] = 3'b110;
        rom_memory[34912] = 3'b110;
        rom_memory[34913] = 3'b110;
        rom_memory[34914] = 3'b110;
        rom_memory[34915] = 3'b110;
        rom_memory[34916] = 3'b110;
        rom_memory[34917] = 3'b110;
        rom_memory[34918] = 3'b110;
        rom_memory[34919] = 3'b110;
        rom_memory[34920] = 3'b110;
        rom_memory[34921] = 3'b110;
        rom_memory[34922] = 3'b110;
        rom_memory[34923] = 3'b110;
        rom_memory[34924] = 3'b110;
        rom_memory[34925] = 3'b110;
        rom_memory[34926] = 3'b110;
        rom_memory[34927] = 3'b110;
        rom_memory[34928] = 3'b110;
        rom_memory[34929] = 3'b110;
        rom_memory[34930] = 3'b110;
        rom_memory[34931] = 3'b110;
        rom_memory[34932] = 3'b110;
        rom_memory[34933] = 3'b110;
        rom_memory[34934] = 3'b110;
        rom_memory[34935] = 3'b110;
        rom_memory[34936] = 3'b110;
        rom_memory[34937] = 3'b110;
        rom_memory[34938] = 3'b110;
        rom_memory[34939] = 3'b110;
        rom_memory[34940] = 3'b110;
        rom_memory[34941] = 3'b110;
        rom_memory[34942] = 3'b110;
        rom_memory[34943] = 3'b110;
        rom_memory[34944] = 3'b110;
        rom_memory[34945] = 3'b000;
        rom_memory[34946] = 3'b000;
        rom_memory[34947] = 3'b000;
        rom_memory[34948] = 3'b000;
        rom_memory[34949] = 3'b000;
        rom_memory[34950] = 3'b110;
        rom_memory[34951] = 3'b110;
        rom_memory[34952] = 3'b000;
        rom_memory[34953] = 3'b000;
        rom_memory[34954] = 3'b110;
        rom_memory[34955] = 3'b100;
        rom_memory[34956] = 3'b000;
        rom_memory[34957] = 3'b000;
        rom_memory[34958] = 3'b100;
        rom_memory[34959] = 3'b110;
        rom_memory[34960] = 3'b111;
        rom_memory[34961] = 3'b110;
        rom_memory[34962] = 3'b110;
        rom_memory[34963] = 3'b110;
        rom_memory[34964] = 3'b110;
        rom_memory[34965] = 3'b110;
        rom_memory[34966] = 3'b110;
        rom_memory[34967] = 3'b110;
        rom_memory[34968] = 3'b110;
        rom_memory[34969] = 3'b110;
        rom_memory[34970] = 3'b110;
        rom_memory[34971] = 3'b110;
        rom_memory[34972] = 3'b110;
        rom_memory[34973] = 3'b110;
        rom_memory[34974] = 3'b110;
        rom_memory[34975] = 3'b110;
        rom_memory[34976] = 3'b110;
        rom_memory[34977] = 3'b110;
        rom_memory[34978] = 3'b110;
        rom_memory[34979] = 3'b110;
        rom_memory[34980] = 3'b110;
        rom_memory[34981] = 3'b110;
        rom_memory[34982] = 3'b110;
        rom_memory[34983] = 3'b110;
        rom_memory[34984] = 3'b110;
        rom_memory[34985] = 3'b110;
        rom_memory[34986] = 3'b110;
        rom_memory[34987] = 3'b110;
        rom_memory[34988] = 3'b111;
        rom_memory[34989] = 3'b110;
        rom_memory[34990] = 3'b110;
        rom_memory[34991] = 3'b110;
        rom_memory[34992] = 3'b110;
        rom_memory[34993] = 3'b111;
        rom_memory[34994] = 3'b111;
        rom_memory[34995] = 3'b111;
        rom_memory[34996] = 3'b111;
        rom_memory[34997] = 3'b111;
        rom_memory[34998] = 3'b111;
        rom_memory[34999] = 3'b111;
        rom_memory[35000] = 3'b111;
        rom_memory[35001] = 3'b111;
        rom_memory[35002] = 3'b111;
        rom_memory[35003] = 3'b111;
        rom_memory[35004] = 3'b111;
        rom_memory[35005] = 3'b111;
        rom_memory[35006] = 3'b111;
        rom_memory[35007] = 3'b111;
        rom_memory[35008] = 3'b111;
        rom_memory[35009] = 3'b111;
        rom_memory[35010] = 3'b111;
        rom_memory[35011] = 3'b111;
        rom_memory[35012] = 3'b111;
        rom_memory[35013] = 3'b111;
        rom_memory[35014] = 3'b111;
        rom_memory[35015] = 3'b111;
        rom_memory[35016] = 3'b111;
        rom_memory[35017] = 3'b111;
        rom_memory[35018] = 3'b111;
        rom_memory[35019] = 3'b111;
        rom_memory[35020] = 3'b111;
        rom_memory[35021] = 3'b111;
        rom_memory[35022] = 3'b111;
        rom_memory[35023] = 3'b111;
        rom_memory[35024] = 3'b111;
        rom_memory[35025] = 3'b111;
        rom_memory[35026] = 3'b111;
        rom_memory[35027] = 3'b111;
        rom_memory[35028] = 3'b111;
        rom_memory[35029] = 3'b111;
        rom_memory[35030] = 3'b111;
        rom_memory[35031] = 3'b111;
        rom_memory[35032] = 3'b111;
        rom_memory[35033] = 3'b111;
        rom_memory[35034] = 3'b111;
        rom_memory[35035] = 3'b111;
        rom_memory[35036] = 3'b111;
        rom_memory[35037] = 3'b111;
        rom_memory[35038] = 3'b111;
        rom_memory[35039] = 3'b111;
        rom_memory[35040] = 3'b110;
        rom_memory[35041] = 3'b110;
        rom_memory[35042] = 3'b110;
        rom_memory[35043] = 3'b110;
        rom_memory[35044] = 3'b110;
        rom_memory[35045] = 3'b111;
        rom_memory[35046] = 3'b111;
        rom_memory[35047] = 3'b111;
        rom_memory[35048] = 3'b111;
        rom_memory[35049] = 3'b111;
        rom_memory[35050] = 3'b111;
        rom_memory[35051] = 3'b111;
        rom_memory[35052] = 3'b111;
        rom_memory[35053] = 3'b111;
        rom_memory[35054] = 3'b111;
        rom_memory[35055] = 3'b111;
        rom_memory[35056] = 3'b111;
        rom_memory[35057] = 3'b111;
        rom_memory[35058] = 3'b111;
        rom_memory[35059] = 3'b111;
        rom_memory[35060] = 3'b111;
        rom_memory[35061] = 3'b111;
        rom_memory[35062] = 3'b111;
        rom_memory[35063] = 3'b110;
        rom_memory[35064] = 3'b110;
        rom_memory[35065] = 3'b110;
        rom_memory[35066] = 3'b110;
        rom_memory[35067] = 3'b110;
        rom_memory[35068] = 3'b111;
        rom_memory[35069] = 3'b111;
        rom_memory[35070] = 3'b111;
        rom_memory[35071] = 3'b110;
        rom_memory[35072] = 3'b110;
        rom_memory[35073] = 3'b110;
        rom_memory[35074] = 3'b110;
        rom_memory[35075] = 3'b110;
        rom_memory[35076] = 3'b110;
        rom_memory[35077] = 3'b110;
        rom_memory[35078] = 3'b110;
        rom_memory[35079] = 3'b110;
        rom_memory[35080] = 3'b110;
        rom_memory[35081] = 3'b110;
        rom_memory[35082] = 3'b110;
        rom_memory[35083] = 3'b110;
        rom_memory[35084] = 3'b111;
        rom_memory[35085] = 3'b111;
        rom_memory[35086] = 3'b111;
        rom_memory[35087] = 3'b111;
        rom_memory[35088] = 3'b111;
        rom_memory[35089] = 3'b111;
        rom_memory[35090] = 3'b111;
        rom_memory[35091] = 3'b111;
        rom_memory[35092] = 3'b111;
        rom_memory[35093] = 3'b111;
        rom_memory[35094] = 3'b111;
        rom_memory[35095] = 3'b110;
        rom_memory[35096] = 3'b111;
        rom_memory[35097] = 3'b111;
        rom_memory[35098] = 3'b111;
        rom_memory[35099] = 3'b111;
        rom_memory[35100] = 3'b111;
        rom_memory[35101] = 3'b111;
        rom_memory[35102] = 3'b111;
        rom_memory[35103] = 3'b000;
        rom_memory[35104] = 3'b000;
        rom_memory[35105] = 3'b000;
        rom_memory[35106] = 3'b000;
        rom_memory[35107] = 3'b000;
        rom_memory[35108] = 3'b000;
        rom_memory[35109] = 3'b000;
        rom_memory[35110] = 3'b000;
        rom_memory[35111] = 3'b000;
        rom_memory[35112] = 3'b000;
        rom_memory[35113] = 3'b000;
        rom_memory[35114] = 3'b000;
        rom_memory[35115] = 3'b111;
        rom_memory[35116] = 3'b100;
        rom_memory[35117] = 3'b000;
        rom_memory[35118] = 3'b110;
        rom_memory[35119] = 3'b100;
        rom_memory[35120] = 3'b100;
        rom_memory[35121] = 3'b100;
        rom_memory[35122] = 3'b111;
        rom_memory[35123] = 3'b000;
        rom_memory[35124] = 3'b000;
        rom_memory[35125] = 3'b000;
        rom_memory[35126] = 3'b000;
        rom_memory[35127] = 3'b110;
        rom_memory[35128] = 3'b100;
        rom_memory[35129] = 3'b111;
        rom_memory[35130] = 3'b111;
        rom_memory[35131] = 3'b111;
        rom_memory[35132] = 3'b111;
        rom_memory[35133] = 3'b111;
        rom_memory[35134] = 3'b110;
        rom_memory[35135] = 3'b110;
        rom_memory[35136] = 3'b110;
        rom_memory[35137] = 3'b111;
        rom_memory[35138] = 3'b110;
        rom_memory[35139] = 3'b110;
        rom_memory[35140] = 3'b110;
        rom_memory[35141] = 3'b110;
        rom_memory[35142] = 3'b110;
        rom_memory[35143] = 3'b110;
        rom_memory[35144] = 3'b110;
        rom_memory[35145] = 3'b110;
        rom_memory[35146] = 3'b110;
        rom_memory[35147] = 3'b110;
        rom_memory[35148] = 3'b110;
        rom_memory[35149] = 3'b110;
        rom_memory[35150] = 3'b110;
        rom_memory[35151] = 3'b110;
        rom_memory[35152] = 3'b110;
        rom_memory[35153] = 3'b110;
        rom_memory[35154] = 3'b110;
        rom_memory[35155] = 3'b110;
        rom_memory[35156] = 3'b110;
        rom_memory[35157] = 3'b110;
        rom_memory[35158] = 3'b110;
        rom_memory[35159] = 3'b110;
        rom_memory[35160] = 3'b110;
        rom_memory[35161] = 3'b110;
        rom_memory[35162] = 3'b110;
        rom_memory[35163] = 3'b110;
        rom_memory[35164] = 3'b110;
        rom_memory[35165] = 3'b110;
        rom_memory[35166] = 3'b110;
        rom_memory[35167] = 3'b110;
        rom_memory[35168] = 3'b110;
        rom_memory[35169] = 3'b110;
        rom_memory[35170] = 3'b110;
        rom_memory[35171] = 3'b110;
        rom_memory[35172] = 3'b110;
        rom_memory[35173] = 3'b110;
        rom_memory[35174] = 3'b110;
        rom_memory[35175] = 3'b110;
        rom_memory[35176] = 3'b110;
        rom_memory[35177] = 3'b110;
        rom_memory[35178] = 3'b110;
        rom_memory[35179] = 3'b110;
        rom_memory[35180] = 3'b110;
        rom_memory[35181] = 3'b110;
        rom_memory[35182] = 3'b110;
        rom_memory[35183] = 3'b110;
        rom_memory[35184] = 3'b110;
        rom_memory[35185] = 3'b110;
        rom_memory[35186] = 3'b000;
        rom_memory[35187] = 3'b000;
        rom_memory[35188] = 3'b000;
        rom_memory[35189] = 3'b000;
        rom_memory[35190] = 3'b000;
        rom_memory[35191] = 3'b110;
        rom_memory[35192] = 3'b110;
        rom_memory[35193] = 3'b000;
        rom_memory[35194] = 3'b000;
        rom_memory[35195] = 3'b110;
        rom_memory[35196] = 3'b000;
        rom_memory[35197] = 3'b000;
        rom_memory[35198] = 3'b000;
        rom_memory[35199] = 3'b000;
        rom_memory[35200] = 3'b110;
        rom_memory[35201] = 3'b110;
        rom_memory[35202] = 3'b110;
        rom_memory[35203] = 3'b110;
        rom_memory[35204] = 3'b110;
        rom_memory[35205] = 3'b110;
        rom_memory[35206] = 3'b110;
        rom_memory[35207] = 3'b110;
        rom_memory[35208] = 3'b110;
        rom_memory[35209] = 3'b110;
        rom_memory[35210] = 3'b110;
        rom_memory[35211] = 3'b110;
        rom_memory[35212] = 3'b110;
        rom_memory[35213] = 3'b110;
        rom_memory[35214] = 3'b110;
        rom_memory[35215] = 3'b110;
        rom_memory[35216] = 3'b110;
        rom_memory[35217] = 3'b110;
        rom_memory[35218] = 3'b110;
        rom_memory[35219] = 3'b110;
        rom_memory[35220] = 3'b110;
        rom_memory[35221] = 3'b110;
        rom_memory[35222] = 3'b110;
        rom_memory[35223] = 3'b110;
        rom_memory[35224] = 3'b110;
        rom_memory[35225] = 3'b110;
        rom_memory[35226] = 3'b110;
        rom_memory[35227] = 3'b110;
        rom_memory[35228] = 3'b110;
        rom_memory[35229] = 3'b110;
        rom_memory[35230] = 3'b110;
        rom_memory[35231] = 3'b110;
        rom_memory[35232] = 3'b110;
        rom_memory[35233] = 3'b111;
        rom_memory[35234] = 3'b110;
        rom_memory[35235] = 3'b111;
        rom_memory[35236] = 3'b111;
        rom_memory[35237] = 3'b111;
        rom_memory[35238] = 3'b111;
        rom_memory[35239] = 3'b111;
        rom_memory[35240] = 3'b111;
        rom_memory[35241] = 3'b111;
        rom_memory[35242] = 3'b111;
        rom_memory[35243] = 3'b111;
        rom_memory[35244] = 3'b111;
        rom_memory[35245] = 3'b111;
        rom_memory[35246] = 3'b111;
        rom_memory[35247] = 3'b111;
        rom_memory[35248] = 3'b111;
        rom_memory[35249] = 3'b111;
        rom_memory[35250] = 3'b111;
        rom_memory[35251] = 3'b111;
        rom_memory[35252] = 3'b111;
        rom_memory[35253] = 3'b111;
        rom_memory[35254] = 3'b111;
        rom_memory[35255] = 3'b111;
        rom_memory[35256] = 3'b111;
        rom_memory[35257] = 3'b111;
        rom_memory[35258] = 3'b111;
        rom_memory[35259] = 3'b111;
        rom_memory[35260] = 3'b111;
        rom_memory[35261] = 3'b111;
        rom_memory[35262] = 3'b111;
        rom_memory[35263] = 3'b111;
        rom_memory[35264] = 3'b111;
        rom_memory[35265] = 3'b111;
        rom_memory[35266] = 3'b111;
        rom_memory[35267] = 3'b111;
        rom_memory[35268] = 3'b111;
        rom_memory[35269] = 3'b111;
        rom_memory[35270] = 3'b111;
        rom_memory[35271] = 3'b111;
        rom_memory[35272] = 3'b111;
        rom_memory[35273] = 3'b111;
        rom_memory[35274] = 3'b111;
        rom_memory[35275] = 3'b111;
        rom_memory[35276] = 3'b111;
        rom_memory[35277] = 3'b111;
        rom_memory[35278] = 3'b111;
        rom_memory[35279] = 3'b111;
        rom_memory[35280] = 3'b110;
        rom_memory[35281] = 3'b110;
        rom_memory[35282] = 3'b110;
        rom_memory[35283] = 3'b110;
        rom_memory[35284] = 3'b110;
        rom_memory[35285] = 3'b110;
        rom_memory[35286] = 3'b111;
        rom_memory[35287] = 3'b111;
        rom_memory[35288] = 3'b111;
        rom_memory[35289] = 3'b111;
        rom_memory[35290] = 3'b111;
        rom_memory[35291] = 3'b111;
        rom_memory[35292] = 3'b111;
        rom_memory[35293] = 3'b111;
        rom_memory[35294] = 3'b111;
        rom_memory[35295] = 3'b111;
        rom_memory[35296] = 3'b111;
        rom_memory[35297] = 3'b111;
        rom_memory[35298] = 3'b111;
        rom_memory[35299] = 3'b111;
        rom_memory[35300] = 3'b111;
        rom_memory[35301] = 3'b111;
        rom_memory[35302] = 3'b111;
        rom_memory[35303] = 3'b110;
        rom_memory[35304] = 3'b110;
        rom_memory[35305] = 3'b110;
        rom_memory[35306] = 3'b110;
        rom_memory[35307] = 3'b110;
        rom_memory[35308] = 3'b111;
        rom_memory[35309] = 3'b110;
        rom_memory[35310] = 3'b110;
        rom_memory[35311] = 3'b110;
        rom_memory[35312] = 3'b110;
        rom_memory[35313] = 3'b110;
        rom_memory[35314] = 3'b110;
        rom_memory[35315] = 3'b110;
        rom_memory[35316] = 3'b110;
        rom_memory[35317] = 3'b110;
        rom_memory[35318] = 3'b110;
        rom_memory[35319] = 3'b110;
        rom_memory[35320] = 3'b110;
        rom_memory[35321] = 3'b110;
        rom_memory[35322] = 3'b110;
        rom_memory[35323] = 3'b110;
        rom_memory[35324] = 3'b111;
        rom_memory[35325] = 3'b111;
        rom_memory[35326] = 3'b111;
        rom_memory[35327] = 3'b111;
        rom_memory[35328] = 3'b111;
        rom_memory[35329] = 3'b111;
        rom_memory[35330] = 3'b111;
        rom_memory[35331] = 3'b111;
        rom_memory[35332] = 3'b111;
        rom_memory[35333] = 3'b111;
        rom_memory[35334] = 3'b111;
        rom_memory[35335] = 3'b111;
        rom_memory[35336] = 3'b111;
        rom_memory[35337] = 3'b111;
        rom_memory[35338] = 3'b111;
        rom_memory[35339] = 3'b111;
        rom_memory[35340] = 3'b111;
        rom_memory[35341] = 3'b111;
        rom_memory[35342] = 3'b111;
        rom_memory[35343] = 3'b000;
        rom_memory[35344] = 3'b000;
        rom_memory[35345] = 3'b000;
        rom_memory[35346] = 3'b000;
        rom_memory[35347] = 3'b000;
        rom_memory[35348] = 3'b000;
        rom_memory[35349] = 3'b000;
        rom_memory[35350] = 3'b000;
        rom_memory[35351] = 3'b000;
        rom_memory[35352] = 3'b000;
        rom_memory[35353] = 3'b000;
        rom_memory[35354] = 3'b000;
        rom_memory[35355] = 3'b111;
        rom_memory[35356] = 3'b111;
        rom_memory[35357] = 3'b000;
        rom_memory[35358] = 3'b100;
        rom_memory[35359] = 3'b110;
        rom_memory[35360] = 3'b100;
        rom_memory[35361] = 3'b000;
        rom_memory[35362] = 3'b111;
        rom_memory[35363] = 3'b000;
        rom_memory[35364] = 3'b000;
        rom_memory[35365] = 3'b000;
        rom_memory[35366] = 3'b100;
        rom_memory[35367] = 3'b100;
        rom_memory[35368] = 3'b000;
        rom_memory[35369] = 3'b110;
        rom_memory[35370] = 3'b111;
        rom_memory[35371] = 3'b111;
        rom_memory[35372] = 3'b111;
        rom_memory[35373] = 3'b110;
        rom_memory[35374] = 3'b100;
        rom_memory[35375] = 3'b110;
        rom_memory[35376] = 3'b110;
        rom_memory[35377] = 3'b110;
        rom_memory[35378] = 3'b110;
        rom_memory[35379] = 3'b110;
        rom_memory[35380] = 3'b110;
        rom_memory[35381] = 3'b110;
        rom_memory[35382] = 3'b110;
        rom_memory[35383] = 3'b110;
        rom_memory[35384] = 3'b110;
        rom_memory[35385] = 3'b110;
        rom_memory[35386] = 3'b110;
        rom_memory[35387] = 3'b110;
        rom_memory[35388] = 3'b110;
        rom_memory[35389] = 3'b110;
        rom_memory[35390] = 3'b110;
        rom_memory[35391] = 3'b110;
        rom_memory[35392] = 3'b110;
        rom_memory[35393] = 3'b110;
        rom_memory[35394] = 3'b110;
        rom_memory[35395] = 3'b110;
        rom_memory[35396] = 3'b110;
        rom_memory[35397] = 3'b110;
        rom_memory[35398] = 3'b110;
        rom_memory[35399] = 3'b110;
        rom_memory[35400] = 3'b110;
        rom_memory[35401] = 3'b110;
        rom_memory[35402] = 3'b110;
        rom_memory[35403] = 3'b110;
        rom_memory[35404] = 3'b110;
        rom_memory[35405] = 3'b110;
        rom_memory[35406] = 3'b110;
        rom_memory[35407] = 3'b110;
        rom_memory[35408] = 3'b110;
        rom_memory[35409] = 3'b110;
        rom_memory[35410] = 3'b110;
        rom_memory[35411] = 3'b110;
        rom_memory[35412] = 3'b110;
        rom_memory[35413] = 3'b110;
        rom_memory[35414] = 3'b110;
        rom_memory[35415] = 3'b110;
        rom_memory[35416] = 3'b110;
        rom_memory[35417] = 3'b110;
        rom_memory[35418] = 3'b110;
        rom_memory[35419] = 3'b110;
        rom_memory[35420] = 3'b110;
        rom_memory[35421] = 3'b110;
        rom_memory[35422] = 3'b110;
        rom_memory[35423] = 3'b110;
        rom_memory[35424] = 3'b110;
        rom_memory[35425] = 3'b110;
        rom_memory[35426] = 3'b110;
        rom_memory[35427] = 3'b000;
        rom_memory[35428] = 3'b000;
        rom_memory[35429] = 3'b000;
        rom_memory[35430] = 3'b000;
        rom_memory[35431] = 3'b000;
        rom_memory[35432] = 3'b110;
        rom_memory[35433] = 3'b110;
        rom_memory[35434] = 3'b000;
        rom_memory[35435] = 3'b000;
        rom_memory[35436] = 3'b110;
        rom_memory[35437] = 3'b000;
        rom_memory[35438] = 3'b000;
        rom_memory[35439] = 3'b000;
        rom_memory[35440] = 3'b000;
        rom_memory[35441] = 3'b110;
        rom_memory[35442] = 3'b110;
        rom_memory[35443] = 3'b110;
        rom_memory[35444] = 3'b110;
        rom_memory[35445] = 3'b110;
        rom_memory[35446] = 3'b110;
        rom_memory[35447] = 3'b110;
        rom_memory[35448] = 3'b110;
        rom_memory[35449] = 3'b110;
        rom_memory[35450] = 3'b110;
        rom_memory[35451] = 3'b110;
        rom_memory[35452] = 3'b110;
        rom_memory[35453] = 3'b110;
        rom_memory[35454] = 3'b110;
        rom_memory[35455] = 3'b110;
        rom_memory[35456] = 3'b110;
        rom_memory[35457] = 3'b110;
        rom_memory[35458] = 3'b110;
        rom_memory[35459] = 3'b110;
        rom_memory[35460] = 3'b110;
        rom_memory[35461] = 3'b110;
        rom_memory[35462] = 3'b110;
        rom_memory[35463] = 3'b110;
        rom_memory[35464] = 3'b110;
        rom_memory[35465] = 3'b110;
        rom_memory[35466] = 3'b110;
        rom_memory[35467] = 3'b110;
        rom_memory[35468] = 3'b110;
        rom_memory[35469] = 3'b110;
        rom_memory[35470] = 3'b110;
        rom_memory[35471] = 3'b110;
        rom_memory[35472] = 3'b110;
        rom_memory[35473] = 3'b110;
        rom_memory[35474] = 3'b110;
        rom_memory[35475] = 3'b110;
        rom_memory[35476] = 3'b110;
        rom_memory[35477] = 3'b111;
        rom_memory[35478] = 3'b111;
        rom_memory[35479] = 3'b111;
        rom_memory[35480] = 3'b111;
        rom_memory[35481] = 3'b111;
        rom_memory[35482] = 3'b111;
        rom_memory[35483] = 3'b111;
        rom_memory[35484] = 3'b111;
        rom_memory[35485] = 3'b111;
        rom_memory[35486] = 3'b111;
        rom_memory[35487] = 3'b111;
        rom_memory[35488] = 3'b111;
        rom_memory[35489] = 3'b111;
        rom_memory[35490] = 3'b111;
        rom_memory[35491] = 3'b111;
        rom_memory[35492] = 3'b111;
        rom_memory[35493] = 3'b111;
        rom_memory[35494] = 3'b111;
        rom_memory[35495] = 3'b111;
        rom_memory[35496] = 3'b111;
        rom_memory[35497] = 3'b111;
        rom_memory[35498] = 3'b111;
        rom_memory[35499] = 3'b111;
        rom_memory[35500] = 3'b111;
        rom_memory[35501] = 3'b111;
        rom_memory[35502] = 3'b111;
        rom_memory[35503] = 3'b111;
        rom_memory[35504] = 3'b111;
        rom_memory[35505] = 3'b111;
        rom_memory[35506] = 3'b111;
        rom_memory[35507] = 3'b111;
        rom_memory[35508] = 3'b111;
        rom_memory[35509] = 3'b111;
        rom_memory[35510] = 3'b111;
        rom_memory[35511] = 3'b111;
        rom_memory[35512] = 3'b111;
        rom_memory[35513] = 3'b111;
        rom_memory[35514] = 3'b111;
        rom_memory[35515] = 3'b111;
        rom_memory[35516] = 3'b111;
        rom_memory[35517] = 3'b111;
        rom_memory[35518] = 3'b111;
        rom_memory[35519] = 3'b111;
        rom_memory[35520] = 3'b110;
        rom_memory[35521] = 3'b110;
        rom_memory[35522] = 3'b110;
        rom_memory[35523] = 3'b110;
        rom_memory[35524] = 3'b110;
        rom_memory[35525] = 3'b110;
        rom_memory[35526] = 3'b111;
        rom_memory[35527] = 3'b111;
        rom_memory[35528] = 3'b111;
        rom_memory[35529] = 3'b111;
        rom_memory[35530] = 3'b111;
        rom_memory[35531] = 3'b111;
        rom_memory[35532] = 3'b111;
        rom_memory[35533] = 3'b111;
        rom_memory[35534] = 3'b111;
        rom_memory[35535] = 3'b111;
        rom_memory[35536] = 3'b111;
        rom_memory[35537] = 3'b111;
        rom_memory[35538] = 3'b111;
        rom_memory[35539] = 3'b111;
        rom_memory[35540] = 3'b111;
        rom_memory[35541] = 3'b111;
        rom_memory[35542] = 3'b110;
        rom_memory[35543] = 3'b110;
        rom_memory[35544] = 3'b110;
        rom_memory[35545] = 3'b110;
        rom_memory[35546] = 3'b110;
        rom_memory[35547] = 3'b110;
        rom_memory[35548] = 3'b110;
        rom_memory[35549] = 3'b110;
        rom_memory[35550] = 3'b110;
        rom_memory[35551] = 3'b110;
        rom_memory[35552] = 3'b110;
        rom_memory[35553] = 3'b110;
        rom_memory[35554] = 3'b110;
        rom_memory[35555] = 3'b110;
        rom_memory[35556] = 3'b110;
        rom_memory[35557] = 3'b110;
        rom_memory[35558] = 3'b110;
        rom_memory[35559] = 3'b110;
        rom_memory[35560] = 3'b110;
        rom_memory[35561] = 3'b110;
        rom_memory[35562] = 3'b110;
        rom_memory[35563] = 3'b111;
        rom_memory[35564] = 3'b111;
        rom_memory[35565] = 3'b111;
        rom_memory[35566] = 3'b110;
        rom_memory[35567] = 3'b111;
        rom_memory[35568] = 3'b111;
        rom_memory[35569] = 3'b111;
        rom_memory[35570] = 3'b111;
        rom_memory[35571] = 3'b111;
        rom_memory[35572] = 3'b111;
        rom_memory[35573] = 3'b111;
        rom_memory[35574] = 3'b111;
        rom_memory[35575] = 3'b000;
        rom_memory[35576] = 3'b111;
        rom_memory[35577] = 3'b111;
        rom_memory[35578] = 3'b110;
        rom_memory[35579] = 3'b111;
        rom_memory[35580] = 3'b111;
        rom_memory[35581] = 3'b110;
        rom_memory[35582] = 3'b110;
        rom_memory[35583] = 3'b000;
        rom_memory[35584] = 3'b000;
        rom_memory[35585] = 3'b000;
        rom_memory[35586] = 3'b000;
        rom_memory[35587] = 3'b000;
        rom_memory[35588] = 3'b000;
        rom_memory[35589] = 3'b111;
        rom_memory[35590] = 3'b101;
        rom_memory[35591] = 3'b000;
        rom_memory[35592] = 3'b000;
        rom_memory[35593] = 3'b000;
        rom_memory[35594] = 3'b111;
        rom_memory[35595] = 3'b111;
        rom_memory[35596] = 3'b111;
        rom_memory[35597] = 3'b111;
        rom_memory[35598] = 3'b000;
        rom_memory[35599] = 3'b000;
        rom_memory[35600] = 3'b111;
        rom_memory[35601] = 3'b000;
        rom_memory[35602] = 3'b101;
        rom_memory[35603] = 3'b000;
        rom_memory[35604] = 3'b000;
        rom_memory[35605] = 3'b000;
        rom_memory[35606] = 3'b000;
        rom_memory[35607] = 3'b100;
        rom_memory[35608] = 3'b100;
        rom_memory[35609] = 3'b111;
        rom_memory[35610] = 3'b111;
        rom_memory[35611] = 3'b111;
        rom_memory[35612] = 3'b111;
        rom_memory[35613] = 3'b111;
        rom_memory[35614] = 3'b111;
        rom_memory[35615] = 3'b111;
        rom_memory[35616] = 3'b110;
        rom_memory[35617] = 3'b110;
        rom_memory[35618] = 3'b110;
        rom_memory[35619] = 3'b110;
        rom_memory[35620] = 3'b110;
        rom_memory[35621] = 3'b110;
        rom_memory[35622] = 3'b110;
        rom_memory[35623] = 3'b110;
        rom_memory[35624] = 3'b110;
        rom_memory[35625] = 3'b110;
        rom_memory[35626] = 3'b110;
        rom_memory[35627] = 3'b110;
        rom_memory[35628] = 3'b110;
        rom_memory[35629] = 3'b110;
        rom_memory[35630] = 3'b110;
        rom_memory[35631] = 3'b110;
        rom_memory[35632] = 3'b110;
        rom_memory[35633] = 3'b110;
        rom_memory[35634] = 3'b110;
        rom_memory[35635] = 3'b110;
        rom_memory[35636] = 3'b110;
        rom_memory[35637] = 3'b110;
        rom_memory[35638] = 3'b110;
        rom_memory[35639] = 3'b110;
        rom_memory[35640] = 3'b110;
        rom_memory[35641] = 3'b110;
        rom_memory[35642] = 3'b110;
        rom_memory[35643] = 3'b110;
        rom_memory[35644] = 3'b110;
        rom_memory[35645] = 3'b110;
        rom_memory[35646] = 3'b110;
        rom_memory[35647] = 3'b110;
        rom_memory[35648] = 3'b110;
        rom_memory[35649] = 3'b110;
        rom_memory[35650] = 3'b110;
        rom_memory[35651] = 3'b110;
        rom_memory[35652] = 3'b110;
        rom_memory[35653] = 3'b110;
        rom_memory[35654] = 3'b110;
        rom_memory[35655] = 3'b110;
        rom_memory[35656] = 3'b110;
        rom_memory[35657] = 3'b110;
        rom_memory[35658] = 3'b110;
        rom_memory[35659] = 3'b110;
        rom_memory[35660] = 3'b110;
        rom_memory[35661] = 3'b110;
        rom_memory[35662] = 3'b110;
        rom_memory[35663] = 3'b110;
        rom_memory[35664] = 3'b110;
        rom_memory[35665] = 3'b110;
        rom_memory[35666] = 3'b110;
        rom_memory[35667] = 3'b110;
        rom_memory[35668] = 3'b000;
        rom_memory[35669] = 3'b000;
        rom_memory[35670] = 3'b000;
        rom_memory[35671] = 3'b000;
        rom_memory[35672] = 3'b000;
        rom_memory[35673] = 3'b111;
        rom_memory[35674] = 3'b111;
        rom_memory[35675] = 3'b000;
        rom_memory[35676] = 3'b000;
        rom_memory[35677] = 3'b110;
        rom_memory[35678] = 3'b000;
        rom_memory[35679] = 3'b000;
        rom_memory[35680] = 3'b000;
        rom_memory[35681] = 3'b000;
        rom_memory[35682] = 3'b110;
        rom_memory[35683] = 3'b111;
        rom_memory[35684] = 3'b110;
        rom_memory[35685] = 3'b110;
        rom_memory[35686] = 3'b110;
        rom_memory[35687] = 3'b110;
        rom_memory[35688] = 3'b110;
        rom_memory[35689] = 3'b110;
        rom_memory[35690] = 3'b110;
        rom_memory[35691] = 3'b110;
        rom_memory[35692] = 3'b110;
        rom_memory[35693] = 3'b110;
        rom_memory[35694] = 3'b110;
        rom_memory[35695] = 3'b110;
        rom_memory[35696] = 3'b110;
        rom_memory[35697] = 3'b110;
        rom_memory[35698] = 3'b110;
        rom_memory[35699] = 3'b110;
        rom_memory[35700] = 3'b110;
        rom_memory[35701] = 3'b110;
        rom_memory[35702] = 3'b110;
        rom_memory[35703] = 3'b110;
        rom_memory[35704] = 3'b110;
        rom_memory[35705] = 3'b110;
        rom_memory[35706] = 3'b110;
        rom_memory[35707] = 3'b110;
        rom_memory[35708] = 3'b110;
        rom_memory[35709] = 3'b110;
        rom_memory[35710] = 3'b110;
        rom_memory[35711] = 3'b110;
        rom_memory[35712] = 3'b110;
        rom_memory[35713] = 3'b110;
        rom_memory[35714] = 3'b110;
        rom_memory[35715] = 3'b110;
        rom_memory[35716] = 3'b111;
        rom_memory[35717] = 3'b111;
        rom_memory[35718] = 3'b111;
        rom_memory[35719] = 3'b111;
        rom_memory[35720] = 3'b111;
        rom_memory[35721] = 3'b111;
        rom_memory[35722] = 3'b111;
        rom_memory[35723] = 3'b111;
        rom_memory[35724] = 3'b111;
        rom_memory[35725] = 3'b111;
        rom_memory[35726] = 3'b111;
        rom_memory[35727] = 3'b111;
        rom_memory[35728] = 3'b111;
        rom_memory[35729] = 3'b111;
        rom_memory[35730] = 3'b111;
        rom_memory[35731] = 3'b111;
        rom_memory[35732] = 3'b111;
        rom_memory[35733] = 3'b111;
        rom_memory[35734] = 3'b111;
        rom_memory[35735] = 3'b111;
        rom_memory[35736] = 3'b111;
        rom_memory[35737] = 3'b111;
        rom_memory[35738] = 3'b111;
        rom_memory[35739] = 3'b111;
        rom_memory[35740] = 3'b111;
        rom_memory[35741] = 3'b111;
        rom_memory[35742] = 3'b111;
        rom_memory[35743] = 3'b111;
        rom_memory[35744] = 3'b111;
        rom_memory[35745] = 3'b111;
        rom_memory[35746] = 3'b111;
        rom_memory[35747] = 3'b111;
        rom_memory[35748] = 3'b111;
        rom_memory[35749] = 3'b111;
        rom_memory[35750] = 3'b111;
        rom_memory[35751] = 3'b111;
        rom_memory[35752] = 3'b111;
        rom_memory[35753] = 3'b111;
        rom_memory[35754] = 3'b111;
        rom_memory[35755] = 3'b111;
        rom_memory[35756] = 3'b111;
        rom_memory[35757] = 3'b111;
        rom_memory[35758] = 3'b111;
        rom_memory[35759] = 3'b111;
        rom_memory[35760] = 3'b110;
        rom_memory[35761] = 3'b110;
        rom_memory[35762] = 3'b110;
        rom_memory[35763] = 3'b110;
        rom_memory[35764] = 3'b110;
        rom_memory[35765] = 3'b110;
        rom_memory[35766] = 3'b111;
        rom_memory[35767] = 3'b111;
        rom_memory[35768] = 3'b111;
        rom_memory[35769] = 3'b111;
        rom_memory[35770] = 3'b111;
        rom_memory[35771] = 3'b111;
        rom_memory[35772] = 3'b111;
        rom_memory[35773] = 3'b111;
        rom_memory[35774] = 3'b111;
        rom_memory[35775] = 3'b111;
        rom_memory[35776] = 3'b111;
        rom_memory[35777] = 3'b111;
        rom_memory[35778] = 3'b111;
        rom_memory[35779] = 3'b111;
        rom_memory[35780] = 3'b111;
        rom_memory[35781] = 3'b111;
        rom_memory[35782] = 3'b110;
        rom_memory[35783] = 3'b110;
        rom_memory[35784] = 3'b110;
        rom_memory[35785] = 3'b110;
        rom_memory[35786] = 3'b110;
        rom_memory[35787] = 3'b110;
        rom_memory[35788] = 3'b110;
        rom_memory[35789] = 3'b110;
        rom_memory[35790] = 3'b110;
        rom_memory[35791] = 3'b110;
        rom_memory[35792] = 3'b110;
        rom_memory[35793] = 3'b110;
        rom_memory[35794] = 3'b110;
        rom_memory[35795] = 3'b110;
        rom_memory[35796] = 3'b110;
        rom_memory[35797] = 3'b110;
        rom_memory[35798] = 3'b110;
        rom_memory[35799] = 3'b110;
        rom_memory[35800] = 3'b110;
        rom_memory[35801] = 3'b110;
        rom_memory[35802] = 3'b110;
        rom_memory[35803] = 3'b110;
        rom_memory[35804] = 3'b111;
        rom_memory[35805] = 3'b111;
        rom_memory[35806] = 3'b111;
        rom_memory[35807] = 3'b111;
        rom_memory[35808] = 3'b111;
        rom_memory[35809] = 3'b111;
        rom_memory[35810] = 3'b111;
        rom_memory[35811] = 3'b111;
        rom_memory[35812] = 3'b111;
        rom_memory[35813] = 3'b111;
        rom_memory[35814] = 3'b111;
        rom_memory[35815] = 3'b000;
        rom_memory[35816] = 3'b111;
        rom_memory[35817] = 3'b110;
        rom_memory[35818] = 3'b110;
        rom_memory[35819] = 3'b110;
        rom_memory[35820] = 3'b111;
        rom_memory[35821] = 3'b110;
        rom_memory[35822] = 3'b110;
        rom_memory[35823] = 3'b000;
        rom_memory[35824] = 3'b000;
        rom_memory[35825] = 3'b000;
        rom_memory[35826] = 3'b000;
        rom_memory[35827] = 3'b000;
        rom_memory[35828] = 3'b000;
        rom_memory[35829] = 3'b100;
        rom_memory[35830] = 3'b000;
        rom_memory[35831] = 3'b000;
        rom_memory[35832] = 3'b000;
        rom_memory[35833] = 3'b000;
        rom_memory[35834] = 3'b111;
        rom_memory[35835] = 3'b111;
        rom_memory[35836] = 3'b111;
        rom_memory[35837] = 3'b111;
        rom_memory[35838] = 3'b000;
        rom_memory[35839] = 3'b000;
        rom_memory[35840] = 3'b100;
        rom_memory[35841] = 3'b100;
        rom_memory[35842] = 3'b000;
        rom_memory[35843] = 3'b100;
        rom_memory[35844] = 3'b111;
        rom_memory[35845] = 3'b000;
        rom_memory[35846] = 3'b000;
        rom_memory[35847] = 3'b111;
        rom_memory[35848] = 3'b100;
        rom_memory[35849] = 3'b110;
        rom_memory[35850] = 3'b111;
        rom_memory[35851] = 3'b111;
        rom_memory[35852] = 3'b111;
        rom_memory[35853] = 3'b111;
        rom_memory[35854] = 3'b111;
        rom_memory[35855] = 3'b110;
        rom_memory[35856] = 3'b110;
        rom_memory[35857] = 3'b110;
        rom_memory[35858] = 3'b110;
        rom_memory[35859] = 3'b110;
        rom_memory[35860] = 3'b110;
        rom_memory[35861] = 3'b110;
        rom_memory[35862] = 3'b110;
        rom_memory[35863] = 3'b110;
        rom_memory[35864] = 3'b110;
        rom_memory[35865] = 3'b110;
        rom_memory[35866] = 3'b110;
        rom_memory[35867] = 3'b110;
        rom_memory[35868] = 3'b110;
        rom_memory[35869] = 3'b110;
        rom_memory[35870] = 3'b110;
        rom_memory[35871] = 3'b110;
        rom_memory[35872] = 3'b110;
        rom_memory[35873] = 3'b110;
        rom_memory[35874] = 3'b110;
        rom_memory[35875] = 3'b110;
        rom_memory[35876] = 3'b110;
        rom_memory[35877] = 3'b110;
        rom_memory[35878] = 3'b110;
        rom_memory[35879] = 3'b110;
        rom_memory[35880] = 3'b110;
        rom_memory[35881] = 3'b110;
        rom_memory[35882] = 3'b110;
        rom_memory[35883] = 3'b110;
        rom_memory[35884] = 3'b110;
        rom_memory[35885] = 3'b110;
        rom_memory[35886] = 3'b110;
        rom_memory[35887] = 3'b110;
        rom_memory[35888] = 3'b110;
        rom_memory[35889] = 3'b110;
        rom_memory[35890] = 3'b110;
        rom_memory[35891] = 3'b110;
        rom_memory[35892] = 3'b110;
        rom_memory[35893] = 3'b110;
        rom_memory[35894] = 3'b110;
        rom_memory[35895] = 3'b110;
        rom_memory[35896] = 3'b110;
        rom_memory[35897] = 3'b110;
        rom_memory[35898] = 3'b110;
        rom_memory[35899] = 3'b110;
        rom_memory[35900] = 3'b110;
        rom_memory[35901] = 3'b110;
        rom_memory[35902] = 3'b110;
        rom_memory[35903] = 3'b110;
        rom_memory[35904] = 3'b110;
        rom_memory[35905] = 3'b110;
        rom_memory[35906] = 3'b110;
        rom_memory[35907] = 3'b110;
        rom_memory[35908] = 3'b110;
        rom_memory[35909] = 3'b000;
        rom_memory[35910] = 3'b000;
        rom_memory[35911] = 3'b000;
        rom_memory[35912] = 3'b000;
        rom_memory[35913] = 3'b000;
        rom_memory[35914] = 3'b110;
        rom_memory[35915] = 3'b111;
        rom_memory[35916] = 3'b000;
        rom_memory[35917] = 3'b000;
        rom_memory[35918] = 3'b110;
        rom_memory[35919] = 3'b000;
        rom_memory[35920] = 3'b000;
        rom_memory[35921] = 3'b000;
        rom_memory[35922] = 3'b000;
        rom_memory[35923] = 3'b110;
        rom_memory[35924] = 3'b110;
        rom_memory[35925] = 3'b110;
        rom_memory[35926] = 3'b110;
        rom_memory[35927] = 3'b110;
        rom_memory[35928] = 3'b110;
        rom_memory[35929] = 3'b110;
        rom_memory[35930] = 3'b110;
        rom_memory[35931] = 3'b110;
        rom_memory[35932] = 3'b110;
        rom_memory[35933] = 3'b110;
        rom_memory[35934] = 3'b110;
        rom_memory[35935] = 3'b110;
        rom_memory[35936] = 3'b110;
        rom_memory[35937] = 3'b110;
        rom_memory[35938] = 3'b110;
        rom_memory[35939] = 3'b110;
        rom_memory[35940] = 3'b110;
        rom_memory[35941] = 3'b110;
        rom_memory[35942] = 3'b110;
        rom_memory[35943] = 3'b110;
        rom_memory[35944] = 3'b110;
        rom_memory[35945] = 3'b110;
        rom_memory[35946] = 3'b110;
        rom_memory[35947] = 3'b110;
        rom_memory[35948] = 3'b110;
        rom_memory[35949] = 3'b110;
        rom_memory[35950] = 3'b110;
        rom_memory[35951] = 3'b110;
        rom_memory[35952] = 3'b110;
        rom_memory[35953] = 3'b110;
        rom_memory[35954] = 3'b110;
        rom_memory[35955] = 3'b111;
        rom_memory[35956] = 3'b111;
        rom_memory[35957] = 3'b111;
        rom_memory[35958] = 3'b111;
        rom_memory[35959] = 3'b111;
        rom_memory[35960] = 3'b111;
        rom_memory[35961] = 3'b111;
        rom_memory[35962] = 3'b111;
        rom_memory[35963] = 3'b111;
        rom_memory[35964] = 3'b111;
        rom_memory[35965] = 3'b111;
        rom_memory[35966] = 3'b111;
        rom_memory[35967] = 3'b111;
        rom_memory[35968] = 3'b111;
        rom_memory[35969] = 3'b111;
        rom_memory[35970] = 3'b111;
        rom_memory[35971] = 3'b111;
        rom_memory[35972] = 3'b111;
        rom_memory[35973] = 3'b111;
        rom_memory[35974] = 3'b111;
        rom_memory[35975] = 3'b111;
        rom_memory[35976] = 3'b111;
        rom_memory[35977] = 3'b111;
        rom_memory[35978] = 3'b111;
        rom_memory[35979] = 3'b111;
        rom_memory[35980] = 3'b111;
        rom_memory[35981] = 3'b111;
        rom_memory[35982] = 3'b111;
        rom_memory[35983] = 3'b111;
        rom_memory[35984] = 3'b111;
        rom_memory[35985] = 3'b111;
        rom_memory[35986] = 3'b111;
        rom_memory[35987] = 3'b111;
        rom_memory[35988] = 3'b111;
        rom_memory[35989] = 3'b111;
        rom_memory[35990] = 3'b111;
        rom_memory[35991] = 3'b111;
        rom_memory[35992] = 3'b111;
        rom_memory[35993] = 3'b111;
        rom_memory[35994] = 3'b111;
        rom_memory[35995] = 3'b111;
        rom_memory[35996] = 3'b111;
        rom_memory[35997] = 3'b111;
        rom_memory[35998] = 3'b111;
        rom_memory[35999] = 3'b111;
        rom_memory[36000] = 3'b110;
        rom_memory[36001] = 3'b110;
        rom_memory[36002] = 3'b110;
        rom_memory[36003] = 3'b110;
        rom_memory[36004] = 3'b110;
        rom_memory[36005] = 3'b110;
        rom_memory[36006] = 3'b111;
        rom_memory[36007] = 3'b111;
        rom_memory[36008] = 3'b111;
        rom_memory[36009] = 3'b111;
        rom_memory[36010] = 3'b111;
        rom_memory[36011] = 3'b111;
        rom_memory[36012] = 3'b111;
        rom_memory[36013] = 3'b111;
        rom_memory[36014] = 3'b111;
        rom_memory[36015] = 3'b111;
        rom_memory[36016] = 3'b111;
        rom_memory[36017] = 3'b111;
        rom_memory[36018] = 3'b111;
        rom_memory[36019] = 3'b111;
        rom_memory[36020] = 3'b111;
        rom_memory[36021] = 3'b111;
        rom_memory[36022] = 3'b111;
        rom_memory[36023] = 3'b110;
        rom_memory[36024] = 3'b110;
        rom_memory[36025] = 3'b110;
        rom_memory[36026] = 3'b110;
        rom_memory[36027] = 3'b110;
        rom_memory[36028] = 3'b110;
        rom_memory[36029] = 3'b110;
        rom_memory[36030] = 3'b110;
        rom_memory[36031] = 3'b110;
        rom_memory[36032] = 3'b110;
        rom_memory[36033] = 3'b110;
        rom_memory[36034] = 3'b110;
        rom_memory[36035] = 3'b110;
        rom_memory[36036] = 3'b110;
        rom_memory[36037] = 3'b110;
        rom_memory[36038] = 3'b110;
        rom_memory[36039] = 3'b110;
        rom_memory[36040] = 3'b110;
        rom_memory[36041] = 3'b110;
        rom_memory[36042] = 3'b110;
        rom_memory[36043] = 3'b110;
        rom_memory[36044] = 3'b110;
        rom_memory[36045] = 3'b111;
        rom_memory[36046] = 3'b111;
        rom_memory[36047] = 3'b111;
        rom_memory[36048] = 3'b111;
        rom_memory[36049] = 3'b111;
        rom_memory[36050] = 3'b111;
        rom_memory[36051] = 3'b111;
        rom_memory[36052] = 3'b111;
        rom_memory[36053] = 3'b111;
        rom_memory[36054] = 3'b111;
        rom_memory[36055] = 3'b000;
        rom_memory[36056] = 3'b110;
        rom_memory[36057] = 3'b110;
        rom_memory[36058] = 3'b110;
        rom_memory[36059] = 3'b110;
        rom_memory[36060] = 3'b110;
        rom_memory[36061] = 3'b110;
        rom_memory[36062] = 3'b111;
        rom_memory[36063] = 3'b110;
        rom_memory[36064] = 3'b000;
        rom_memory[36065] = 3'b000;
        rom_memory[36066] = 3'b000;
        rom_memory[36067] = 3'b000;
        rom_memory[36068] = 3'b000;
        rom_memory[36069] = 3'b000;
        rom_memory[36070] = 3'b000;
        rom_memory[36071] = 3'b111;
        rom_memory[36072] = 3'b000;
        rom_memory[36073] = 3'b100;
        rom_memory[36074] = 3'b111;
        rom_memory[36075] = 3'b111;
        rom_memory[36076] = 3'b111;
        rom_memory[36077] = 3'b111;
        rom_memory[36078] = 3'b111;
        rom_memory[36079] = 3'b110;
        rom_memory[36080] = 3'b000;
        rom_memory[36081] = 3'b000;
        rom_memory[36082] = 3'b000;
        rom_memory[36083] = 3'b100;
        rom_memory[36084] = 3'b110;
        rom_memory[36085] = 3'b000;
        rom_memory[36086] = 3'b000;
        rom_memory[36087] = 3'b000;
        rom_memory[36088] = 3'b000;
        rom_memory[36089] = 3'b000;
        rom_memory[36090] = 3'b110;
        rom_memory[36091] = 3'b111;
        rom_memory[36092] = 3'b111;
        rom_memory[36093] = 3'b111;
        rom_memory[36094] = 3'b110;
        rom_memory[36095] = 3'b110;
        rom_memory[36096] = 3'b110;
        rom_memory[36097] = 3'b110;
        rom_memory[36098] = 3'b110;
        rom_memory[36099] = 3'b110;
        rom_memory[36100] = 3'b110;
        rom_memory[36101] = 3'b110;
        rom_memory[36102] = 3'b110;
        rom_memory[36103] = 3'b110;
        rom_memory[36104] = 3'b110;
        rom_memory[36105] = 3'b110;
        rom_memory[36106] = 3'b110;
        rom_memory[36107] = 3'b110;
        rom_memory[36108] = 3'b110;
        rom_memory[36109] = 3'b110;
        rom_memory[36110] = 3'b110;
        rom_memory[36111] = 3'b110;
        rom_memory[36112] = 3'b110;
        rom_memory[36113] = 3'b110;
        rom_memory[36114] = 3'b110;
        rom_memory[36115] = 3'b110;
        rom_memory[36116] = 3'b110;
        rom_memory[36117] = 3'b110;
        rom_memory[36118] = 3'b110;
        rom_memory[36119] = 3'b110;
        rom_memory[36120] = 3'b110;
        rom_memory[36121] = 3'b110;
        rom_memory[36122] = 3'b110;
        rom_memory[36123] = 3'b110;
        rom_memory[36124] = 3'b110;
        rom_memory[36125] = 3'b110;
        rom_memory[36126] = 3'b110;
        rom_memory[36127] = 3'b110;
        rom_memory[36128] = 3'b110;
        rom_memory[36129] = 3'b110;
        rom_memory[36130] = 3'b110;
        rom_memory[36131] = 3'b110;
        rom_memory[36132] = 3'b110;
        rom_memory[36133] = 3'b110;
        rom_memory[36134] = 3'b110;
        rom_memory[36135] = 3'b110;
        rom_memory[36136] = 3'b110;
        rom_memory[36137] = 3'b110;
        rom_memory[36138] = 3'b110;
        rom_memory[36139] = 3'b110;
        rom_memory[36140] = 3'b110;
        rom_memory[36141] = 3'b110;
        rom_memory[36142] = 3'b110;
        rom_memory[36143] = 3'b110;
        rom_memory[36144] = 3'b110;
        rom_memory[36145] = 3'b110;
        rom_memory[36146] = 3'b110;
        rom_memory[36147] = 3'b110;
        rom_memory[36148] = 3'b110;
        rom_memory[36149] = 3'b110;
        rom_memory[36150] = 3'b000;
        rom_memory[36151] = 3'b000;
        rom_memory[36152] = 3'b000;
        rom_memory[36153] = 3'b000;
        rom_memory[36154] = 3'b000;
        rom_memory[36155] = 3'b110;
        rom_memory[36156] = 3'b111;
        rom_memory[36157] = 3'b000;
        rom_memory[36158] = 3'b000;
        rom_memory[36159] = 3'b110;
        rom_memory[36160] = 3'b000;
        rom_memory[36161] = 3'b000;
        rom_memory[36162] = 3'b000;
        rom_memory[36163] = 3'b000;
        rom_memory[36164] = 3'b110;
        rom_memory[36165] = 3'b111;
        rom_memory[36166] = 3'b110;
        rom_memory[36167] = 3'b110;
        rom_memory[36168] = 3'b110;
        rom_memory[36169] = 3'b110;
        rom_memory[36170] = 3'b110;
        rom_memory[36171] = 3'b110;
        rom_memory[36172] = 3'b110;
        rom_memory[36173] = 3'b110;
        rom_memory[36174] = 3'b110;
        rom_memory[36175] = 3'b110;
        rom_memory[36176] = 3'b110;
        rom_memory[36177] = 3'b110;
        rom_memory[36178] = 3'b110;
        rom_memory[36179] = 3'b110;
        rom_memory[36180] = 3'b110;
        rom_memory[36181] = 3'b110;
        rom_memory[36182] = 3'b110;
        rom_memory[36183] = 3'b110;
        rom_memory[36184] = 3'b110;
        rom_memory[36185] = 3'b110;
        rom_memory[36186] = 3'b110;
        rom_memory[36187] = 3'b110;
        rom_memory[36188] = 3'b110;
        rom_memory[36189] = 3'b110;
        rom_memory[36190] = 3'b110;
        rom_memory[36191] = 3'b110;
        rom_memory[36192] = 3'b110;
        rom_memory[36193] = 3'b110;
        rom_memory[36194] = 3'b110;
        rom_memory[36195] = 3'b111;
        rom_memory[36196] = 3'b111;
        rom_memory[36197] = 3'b111;
        rom_memory[36198] = 3'b111;
        rom_memory[36199] = 3'b111;
        rom_memory[36200] = 3'b111;
        rom_memory[36201] = 3'b111;
        rom_memory[36202] = 3'b111;
        rom_memory[36203] = 3'b111;
        rom_memory[36204] = 3'b111;
        rom_memory[36205] = 3'b111;
        rom_memory[36206] = 3'b111;
        rom_memory[36207] = 3'b111;
        rom_memory[36208] = 3'b111;
        rom_memory[36209] = 3'b111;
        rom_memory[36210] = 3'b111;
        rom_memory[36211] = 3'b111;
        rom_memory[36212] = 3'b111;
        rom_memory[36213] = 3'b111;
        rom_memory[36214] = 3'b111;
        rom_memory[36215] = 3'b111;
        rom_memory[36216] = 3'b111;
        rom_memory[36217] = 3'b111;
        rom_memory[36218] = 3'b111;
        rom_memory[36219] = 3'b111;
        rom_memory[36220] = 3'b111;
        rom_memory[36221] = 3'b111;
        rom_memory[36222] = 3'b111;
        rom_memory[36223] = 3'b111;
        rom_memory[36224] = 3'b111;
        rom_memory[36225] = 3'b111;
        rom_memory[36226] = 3'b111;
        rom_memory[36227] = 3'b111;
        rom_memory[36228] = 3'b111;
        rom_memory[36229] = 3'b111;
        rom_memory[36230] = 3'b111;
        rom_memory[36231] = 3'b111;
        rom_memory[36232] = 3'b111;
        rom_memory[36233] = 3'b111;
        rom_memory[36234] = 3'b111;
        rom_memory[36235] = 3'b111;
        rom_memory[36236] = 3'b111;
        rom_memory[36237] = 3'b111;
        rom_memory[36238] = 3'b111;
        rom_memory[36239] = 3'b111;
        rom_memory[36240] = 3'b110;
        rom_memory[36241] = 3'b110;
        rom_memory[36242] = 3'b110;
        rom_memory[36243] = 3'b110;
        rom_memory[36244] = 3'b110;
        rom_memory[36245] = 3'b110;
        rom_memory[36246] = 3'b111;
        rom_memory[36247] = 3'b111;
        rom_memory[36248] = 3'b111;
        rom_memory[36249] = 3'b111;
        rom_memory[36250] = 3'b111;
        rom_memory[36251] = 3'b111;
        rom_memory[36252] = 3'b111;
        rom_memory[36253] = 3'b111;
        rom_memory[36254] = 3'b111;
        rom_memory[36255] = 3'b111;
        rom_memory[36256] = 3'b111;
        rom_memory[36257] = 3'b111;
        rom_memory[36258] = 3'b111;
        rom_memory[36259] = 3'b111;
        rom_memory[36260] = 3'b111;
        rom_memory[36261] = 3'b111;
        rom_memory[36262] = 3'b111;
        rom_memory[36263] = 3'b110;
        rom_memory[36264] = 3'b110;
        rom_memory[36265] = 3'b110;
        rom_memory[36266] = 3'b110;
        rom_memory[36267] = 3'b110;
        rom_memory[36268] = 3'b110;
        rom_memory[36269] = 3'b110;
        rom_memory[36270] = 3'b110;
        rom_memory[36271] = 3'b110;
        rom_memory[36272] = 3'b110;
        rom_memory[36273] = 3'b110;
        rom_memory[36274] = 3'b110;
        rom_memory[36275] = 3'b110;
        rom_memory[36276] = 3'b110;
        rom_memory[36277] = 3'b110;
        rom_memory[36278] = 3'b110;
        rom_memory[36279] = 3'b110;
        rom_memory[36280] = 3'b110;
        rom_memory[36281] = 3'b110;
        rom_memory[36282] = 3'b110;
        rom_memory[36283] = 3'b111;
        rom_memory[36284] = 3'b111;
        rom_memory[36285] = 3'b111;
        rom_memory[36286] = 3'b110;
        rom_memory[36287] = 3'b110;
        rom_memory[36288] = 3'b110;
        rom_memory[36289] = 3'b111;
        rom_memory[36290] = 3'b111;
        rom_memory[36291] = 3'b111;
        rom_memory[36292] = 3'b111;
        rom_memory[36293] = 3'b111;
        rom_memory[36294] = 3'b111;
        rom_memory[36295] = 3'b000;
        rom_memory[36296] = 3'b110;
        rom_memory[36297] = 3'b110;
        rom_memory[36298] = 3'b110;
        rom_memory[36299] = 3'b110;
        rom_memory[36300] = 3'b110;
        rom_memory[36301] = 3'b111;
        rom_memory[36302] = 3'b111;
        rom_memory[36303] = 3'b110;
        rom_memory[36304] = 3'b111;
        rom_memory[36305] = 3'b111;
        rom_memory[36306] = 3'b000;
        rom_memory[36307] = 3'b000;
        rom_memory[36308] = 3'b100;
        rom_memory[36309] = 3'b110;
        rom_memory[36310] = 3'b111;
        rom_memory[36311] = 3'b100;
        rom_memory[36312] = 3'b000;
        rom_memory[36313] = 3'b110;
        rom_memory[36314] = 3'b111;
        rom_memory[36315] = 3'b111;
        rom_memory[36316] = 3'b110;
        rom_memory[36317] = 3'b110;
        rom_memory[36318] = 3'b110;
        rom_memory[36319] = 3'b110;
        rom_memory[36320] = 3'b000;
        rom_memory[36321] = 3'b000;
        rom_memory[36322] = 3'b000;
        rom_memory[36323] = 3'b000;
        rom_memory[36324] = 3'b000;
        rom_memory[36325] = 3'b000;
        rom_memory[36326] = 3'b000;
        rom_memory[36327] = 3'b000;
        rom_memory[36328] = 3'b000;
        rom_memory[36329] = 3'b000;
        rom_memory[36330] = 3'b100;
        rom_memory[36331] = 3'b111;
        rom_memory[36332] = 3'b000;
        rom_memory[36333] = 3'b000;
        rom_memory[36334] = 3'b000;
        rom_memory[36335] = 3'b110;
        rom_memory[36336] = 3'b110;
        rom_memory[36337] = 3'b110;
        rom_memory[36338] = 3'b110;
        rom_memory[36339] = 3'b110;
        rom_memory[36340] = 3'b110;
        rom_memory[36341] = 3'b110;
        rom_memory[36342] = 3'b110;
        rom_memory[36343] = 3'b110;
        rom_memory[36344] = 3'b110;
        rom_memory[36345] = 3'b110;
        rom_memory[36346] = 3'b110;
        rom_memory[36347] = 3'b110;
        rom_memory[36348] = 3'b110;
        rom_memory[36349] = 3'b110;
        rom_memory[36350] = 3'b110;
        rom_memory[36351] = 3'b110;
        rom_memory[36352] = 3'b110;
        rom_memory[36353] = 3'b110;
        rom_memory[36354] = 3'b110;
        rom_memory[36355] = 3'b110;
        rom_memory[36356] = 3'b110;
        rom_memory[36357] = 3'b110;
        rom_memory[36358] = 3'b110;
        rom_memory[36359] = 3'b110;
        rom_memory[36360] = 3'b110;
        rom_memory[36361] = 3'b110;
        rom_memory[36362] = 3'b110;
        rom_memory[36363] = 3'b110;
        rom_memory[36364] = 3'b110;
        rom_memory[36365] = 3'b110;
        rom_memory[36366] = 3'b110;
        rom_memory[36367] = 3'b110;
        rom_memory[36368] = 3'b110;
        rom_memory[36369] = 3'b110;
        rom_memory[36370] = 3'b110;
        rom_memory[36371] = 3'b110;
        rom_memory[36372] = 3'b110;
        rom_memory[36373] = 3'b110;
        rom_memory[36374] = 3'b110;
        rom_memory[36375] = 3'b110;
        rom_memory[36376] = 3'b110;
        rom_memory[36377] = 3'b110;
        rom_memory[36378] = 3'b110;
        rom_memory[36379] = 3'b110;
        rom_memory[36380] = 3'b110;
        rom_memory[36381] = 3'b110;
        rom_memory[36382] = 3'b110;
        rom_memory[36383] = 3'b110;
        rom_memory[36384] = 3'b110;
        rom_memory[36385] = 3'b110;
        rom_memory[36386] = 3'b110;
        rom_memory[36387] = 3'b110;
        rom_memory[36388] = 3'b110;
        rom_memory[36389] = 3'b110;
        rom_memory[36390] = 3'b110;
        rom_memory[36391] = 3'b000;
        rom_memory[36392] = 3'b000;
        rom_memory[36393] = 3'b000;
        rom_memory[36394] = 3'b000;
        rom_memory[36395] = 3'b000;
        rom_memory[36396] = 3'b110;
        rom_memory[36397] = 3'b111;
        rom_memory[36398] = 3'b000;
        rom_memory[36399] = 3'b000;
        rom_memory[36400] = 3'b110;
        rom_memory[36401] = 3'b000;
        rom_memory[36402] = 3'b000;
        rom_memory[36403] = 3'b000;
        rom_memory[36404] = 3'b000;
        rom_memory[36405] = 3'b110;
        rom_memory[36406] = 3'b111;
        rom_memory[36407] = 3'b110;
        rom_memory[36408] = 3'b110;
        rom_memory[36409] = 3'b110;
        rom_memory[36410] = 3'b110;
        rom_memory[36411] = 3'b110;
        rom_memory[36412] = 3'b110;
        rom_memory[36413] = 3'b110;
        rom_memory[36414] = 3'b110;
        rom_memory[36415] = 3'b110;
        rom_memory[36416] = 3'b110;
        rom_memory[36417] = 3'b110;
        rom_memory[36418] = 3'b110;
        rom_memory[36419] = 3'b110;
        rom_memory[36420] = 3'b110;
        rom_memory[36421] = 3'b110;
        rom_memory[36422] = 3'b110;
        rom_memory[36423] = 3'b110;
        rom_memory[36424] = 3'b110;
        rom_memory[36425] = 3'b110;
        rom_memory[36426] = 3'b110;
        rom_memory[36427] = 3'b110;
        rom_memory[36428] = 3'b110;
        rom_memory[36429] = 3'b110;
        rom_memory[36430] = 3'b110;
        rom_memory[36431] = 3'b110;
        rom_memory[36432] = 3'b110;
        rom_memory[36433] = 3'b110;
        rom_memory[36434] = 3'b110;
        rom_memory[36435] = 3'b111;
        rom_memory[36436] = 3'b111;
        rom_memory[36437] = 3'b111;
        rom_memory[36438] = 3'b110;
        rom_memory[36439] = 3'b111;
        rom_memory[36440] = 3'b111;
        rom_memory[36441] = 3'b111;
        rom_memory[36442] = 3'b111;
        rom_memory[36443] = 3'b111;
        rom_memory[36444] = 3'b111;
        rom_memory[36445] = 3'b111;
        rom_memory[36446] = 3'b111;
        rom_memory[36447] = 3'b111;
        rom_memory[36448] = 3'b111;
        rom_memory[36449] = 3'b111;
        rom_memory[36450] = 3'b111;
        rom_memory[36451] = 3'b111;
        rom_memory[36452] = 3'b111;
        rom_memory[36453] = 3'b111;
        rom_memory[36454] = 3'b111;
        rom_memory[36455] = 3'b111;
        rom_memory[36456] = 3'b111;
        rom_memory[36457] = 3'b111;
        rom_memory[36458] = 3'b111;
        rom_memory[36459] = 3'b111;
        rom_memory[36460] = 3'b111;
        rom_memory[36461] = 3'b111;
        rom_memory[36462] = 3'b111;
        rom_memory[36463] = 3'b111;
        rom_memory[36464] = 3'b111;
        rom_memory[36465] = 3'b111;
        rom_memory[36466] = 3'b111;
        rom_memory[36467] = 3'b111;
        rom_memory[36468] = 3'b111;
        rom_memory[36469] = 3'b111;
        rom_memory[36470] = 3'b111;
        rom_memory[36471] = 3'b111;
        rom_memory[36472] = 3'b111;
        rom_memory[36473] = 3'b111;
        rom_memory[36474] = 3'b111;
        rom_memory[36475] = 3'b111;
        rom_memory[36476] = 3'b111;
        rom_memory[36477] = 3'b111;
        rom_memory[36478] = 3'b111;
        rom_memory[36479] = 3'b111;
        rom_memory[36480] = 3'b110;
        rom_memory[36481] = 3'b110;
        rom_memory[36482] = 3'b110;
        rom_memory[36483] = 3'b110;
        rom_memory[36484] = 3'b110;
        rom_memory[36485] = 3'b110;
        rom_memory[36486] = 3'b111;
        rom_memory[36487] = 3'b111;
        rom_memory[36488] = 3'b111;
        rom_memory[36489] = 3'b111;
        rom_memory[36490] = 3'b111;
        rom_memory[36491] = 3'b111;
        rom_memory[36492] = 3'b111;
        rom_memory[36493] = 3'b111;
        rom_memory[36494] = 3'b111;
        rom_memory[36495] = 3'b111;
        rom_memory[36496] = 3'b111;
        rom_memory[36497] = 3'b111;
        rom_memory[36498] = 3'b111;
        rom_memory[36499] = 3'b111;
        rom_memory[36500] = 3'b111;
        rom_memory[36501] = 3'b111;
        rom_memory[36502] = 3'b111;
        rom_memory[36503] = 3'b111;
        rom_memory[36504] = 3'b110;
        rom_memory[36505] = 3'b110;
        rom_memory[36506] = 3'b110;
        rom_memory[36507] = 3'b110;
        rom_memory[36508] = 3'b110;
        rom_memory[36509] = 3'b110;
        rom_memory[36510] = 3'b110;
        rom_memory[36511] = 3'b110;
        rom_memory[36512] = 3'b110;
        rom_memory[36513] = 3'b110;
        rom_memory[36514] = 3'b110;
        rom_memory[36515] = 3'b110;
        rom_memory[36516] = 3'b110;
        rom_memory[36517] = 3'b110;
        rom_memory[36518] = 3'b110;
        rom_memory[36519] = 3'b110;
        rom_memory[36520] = 3'b110;
        rom_memory[36521] = 3'b110;
        rom_memory[36522] = 3'b110;
        rom_memory[36523] = 3'b110;
        rom_memory[36524] = 3'b111;
        rom_memory[36525] = 3'b111;
        rom_memory[36526] = 3'b111;
        rom_memory[36527] = 3'b111;
        rom_memory[36528] = 3'b110;
        rom_memory[36529] = 3'b110;
        rom_memory[36530] = 3'b110;
        rom_memory[36531] = 3'b110;
        rom_memory[36532] = 3'b110;
        rom_memory[36533] = 3'b111;
        rom_memory[36534] = 3'b111;
        rom_memory[36535] = 3'b000;
        rom_memory[36536] = 3'b110;
        rom_memory[36537] = 3'b110;
        rom_memory[36538] = 3'b110;
        rom_memory[36539] = 3'b110;
        rom_memory[36540] = 3'b110;
        rom_memory[36541] = 3'b111;
        rom_memory[36542] = 3'b111;
        rom_memory[36543] = 3'b110;
        rom_memory[36544] = 3'b111;
        rom_memory[36545] = 3'b110;
        rom_memory[36546] = 3'b000;
        rom_memory[36547] = 3'b000;
        rom_memory[36548] = 3'b000;
        rom_memory[36549] = 3'b111;
        rom_memory[36550] = 3'b110;
        rom_memory[36551] = 3'b110;
        rom_memory[36552] = 3'b110;
        rom_memory[36553] = 3'b111;
        rom_memory[36554] = 3'b111;
        rom_memory[36555] = 3'b111;
        rom_memory[36556] = 3'b111;
        rom_memory[36557] = 3'b110;
        rom_memory[36558] = 3'b110;
        rom_memory[36559] = 3'b110;
        rom_memory[36560] = 3'b100;
        rom_memory[36561] = 3'b000;
        rom_memory[36562] = 3'b000;
        rom_memory[36563] = 3'b000;
        rom_memory[36564] = 3'b000;
        rom_memory[36565] = 3'b000;
        rom_memory[36566] = 3'b000;
        rom_memory[36567] = 3'b000;
        rom_memory[36568] = 3'b111;
        rom_memory[36569] = 3'b000;
        rom_memory[36570] = 3'b100;
        rom_memory[36571] = 3'b111;
        rom_memory[36572] = 3'b101;
        rom_memory[36573] = 3'b000;
        rom_memory[36574] = 3'b000;
        rom_memory[36575] = 3'b110;
        rom_memory[36576] = 3'b110;
        rom_memory[36577] = 3'b110;
        rom_memory[36578] = 3'b110;
        rom_memory[36579] = 3'b110;
        rom_memory[36580] = 3'b110;
        rom_memory[36581] = 3'b110;
        rom_memory[36582] = 3'b110;
        rom_memory[36583] = 3'b110;
        rom_memory[36584] = 3'b110;
        rom_memory[36585] = 3'b110;
        rom_memory[36586] = 3'b110;
        rom_memory[36587] = 3'b110;
        rom_memory[36588] = 3'b110;
        rom_memory[36589] = 3'b110;
        rom_memory[36590] = 3'b110;
        rom_memory[36591] = 3'b110;
        rom_memory[36592] = 3'b110;
        rom_memory[36593] = 3'b110;
        rom_memory[36594] = 3'b110;
        rom_memory[36595] = 3'b110;
        rom_memory[36596] = 3'b110;
        rom_memory[36597] = 3'b110;
        rom_memory[36598] = 3'b110;
        rom_memory[36599] = 3'b110;
        rom_memory[36600] = 3'b110;
        rom_memory[36601] = 3'b110;
        rom_memory[36602] = 3'b110;
        rom_memory[36603] = 3'b110;
        rom_memory[36604] = 3'b110;
        rom_memory[36605] = 3'b110;
        rom_memory[36606] = 3'b110;
        rom_memory[36607] = 3'b110;
        rom_memory[36608] = 3'b110;
        rom_memory[36609] = 3'b110;
        rom_memory[36610] = 3'b110;
        rom_memory[36611] = 3'b110;
        rom_memory[36612] = 3'b110;
        rom_memory[36613] = 3'b110;
        rom_memory[36614] = 3'b110;
        rom_memory[36615] = 3'b110;
        rom_memory[36616] = 3'b110;
        rom_memory[36617] = 3'b110;
        rom_memory[36618] = 3'b110;
        rom_memory[36619] = 3'b110;
        rom_memory[36620] = 3'b110;
        rom_memory[36621] = 3'b110;
        rom_memory[36622] = 3'b110;
        rom_memory[36623] = 3'b110;
        rom_memory[36624] = 3'b110;
        rom_memory[36625] = 3'b110;
        rom_memory[36626] = 3'b110;
        rom_memory[36627] = 3'b110;
        rom_memory[36628] = 3'b110;
        rom_memory[36629] = 3'b110;
        rom_memory[36630] = 3'b110;
        rom_memory[36631] = 3'b110;
        rom_memory[36632] = 3'b000;
        rom_memory[36633] = 3'b000;
        rom_memory[36634] = 3'b000;
        rom_memory[36635] = 3'b000;
        rom_memory[36636] = 3'b000;
        rom_memory[36637] = 3'b110;
        rom_memory[36638] = 3'b111;
        rom_memory[36639] = 3'b000;
        rom_memory[36640] = 3'b000;
        rom_memory[36641] = 3'b110;
        rom_memory[36642] = 3'b000;
        rom_memory[36643] = 3'b000;
        rom_memory[36644] = 3'b000;
        rom_memory[36645] = 3'b000;
        rom_memory[36646] = 3'b110;
        rom_memory[36647] = 3'b111;
        rom_memory[36648] = 3'b111;
        rom_memory[36649] = 3'b110;
        rom_memory[36650] = 3'b110;
        rom_memory[36651] = 3'b110;
        rom_memory[36652] = 3'b110;
        rom_memory[36653] = 3'b110;
        rom_memory[36654] = 3'b110;
        rom_memory[36655] = 3'b110;
        rom_memory[36656] = 3'b110;
        rom_memory[36657] = 3'b110;
        rom_memory[36658] = 3'b110;
        rom_memory[36659] = 3'b110;
        rom_memory[36660] = 3'b110;
        rom_memory[36661] = 3'b110;
        rom_memory[36662] = 3'b110;
        rom_memory[36663] = 3'b110;
        rom_memory[36664] = 3'b110;
        rom_memory[36665] = 3'b110;
        rom_memory[36666] = 3'b110;
        rom_memory[36667] = 3'b110;
        rom_memory[36668] = 3'b110;
        rom_memory[36669] = 3'b110;
        rom_memory[36670] = 3'b110;
        rom_memory[36671] = 3'b110;
        rom_memory[36672] = 3'b110;
        rom_memory[36673] = 3'b110;
        rom_memory[36674] = 3'b110;
        rom_memory[36675] = 3'b110;
        rom_memory[36676] = 3'b110;
        rom_memory[36677] = 3'b110;
        rom_memory[36678] = 3'b111;
        rom_memory[36679] = 3'b111;
        rom_memory[36680] = 3'b111;
        rom_memory[36681] = 3'b111;
        rom_memory[36682] = 3'b111;
        rom_memory[36683] = 3'b111;
        rom_memory[36684] = 3'b111;
        rom_memory[36685] = 3'b111;
        rom_memory[36686] = 3'b111;
        rom_memory[36687] = 3'b111;
        rom_memory[36688] = 3'b111;
        rom_memory[36689] = 3'b111;
        rom_memory[36690] = 3'b111;
        rom_memory[36691] = 3'b111;
        rom_memory[36692] = 3'b111;
        rom_memory[36693] = 3'b111;
        rom_memory[36694] = 3'b111;
        rom_memory[36695] = 3'b111;
        rom_memory[36696] = 3'b111;
        rom_memory[36697] = 3'b111;
        rom_memory[36698] = 3'b111;
        rom_memory[36699] = 3'b111;
        rom_memory[36700] = 3'b111;
        rom_memory[36701] = 3'b111;
        rom_memory[36702] = 3'b111;
        rom_memory[36703] = 3'b111;
        rom_memory[36704] = 3'b111;
        rom_memory[36705] = 3'b111;
        rom_memory[36706] = 3'b111;
        rom_memory[36707] = 3'b111;
        rom_memory[36708] = 3'b111;
        rom_memory[36709] = 3'b111;
        rom_memory[36710] = 3'b111;
        rom_memory[36711] = 3'b111;
        rom_memory[36712] = 3'b111;
        rom_memory[36713] = 3'b111;
        rom_memory[36714] = 3'b111;
        rom_memory[36715] = 3'b111;
        rom_memory[36716] = 3'b111;
        rom_memory[36717] = 3'b111;
        rom_memory[36718] = 3'b111;
        rom_memory[36719] = 3'b111;
        rom_memory[36720] = 3'b110;
        rom_memory[36721] = 3'b110;
        rom_memory[36722] = 3'b110;
        rom_memory[36723] = 3'b110;
        rom_memory[36724] = 3'b110;
        rom_memory[36725] = 3'b110;
        rom_memory[36726] = 3'b111;
        rom_memory[36727] = 3'b111;
        rom_memory[36728] = 3'b111;
        rom_memory[36729] = 3'b111;
        rom_memory[36730] = 3'b111;
        rom_memory[36731] = 3'b111;
        rom_memory[36732] = 3'b111;
        rom_memory[36733] = 3'b111;
        rom_memory[36734] = 3'b111;
        rom_memory[36735] = 3'b111;
        rom_memory[36736] = 3'b111;
        rom_memory[36737] = 3'b111;
        rom_memory[36738] = 3'b111;
        rom_memory[36739] = 3'b111;
        rom_memory[36740] = 3'b111;
        rom_memory[36741] = 3'b111;
        rom_memory[36742] = 3'b111;
        rom_memory[36743] = 3'b111;
        rom_memory[36744] = 3'b110;
        rom_memory[36745] = 3'b110;
        rom_memory[36746] = 3'b110;
        rom_memory[36747] = 3'b110;
        rom_memory[36748] = 3'b110;
        rom_memory[36749] = 3'b110;
        rom_memory[36750] = 3'b110;
        rom_memory[36751] = 3'b110;
        rom_memory[36752] = 3'b110;
        rom_memory[36753] = 3'b110;
        rom_memory[36754] = 3'b110;
        rom_memory[36755] = 3'b110;
        rom_memory[36756] = 3'b110;
        rom_memory[36757] = 3'b110;
        rom_memory[36758] = 3'b110;
        rom_memory[36759] = 3'b110;
        rom_memory[36760] = 3'b110;
        rom_memory[36761] = 3'b110;
        rom_memory[36762] = 3'b110;
        rom_memory[36763] = 3'b110;
        rom_memory[36764] = 3'b111;
        rom_memory[36765] = 3'b111;
        rom_memory[36766] = 3'b111;
        rom_memory[36767] = 3'b111;
        rom_memory[36768] = 3'b111;
        rom_memory[36769] = 3'b111;
        rom_memory[36770] = 3'b110;
        rom_memory[36771] = 3'b110;
        rom_memory[36772] = 3'b110;
        rom_memory[36773] = 3'b110;
        rom_memory[36774] = 3'b110;
        rom_memory[36775] = 3'b000;
        rom_memory[36776] = 3'b000;
        rom_memory[36777] = 3'b111;
        rom_memory[36778] = 3'b110;
        rom_memory[36779] = 3'b110;
        rom_memory[36780] = 3'b110;
        rom_memory[36781] = 3'b111;
        rom_memory[36782] = 3'b111;
        rom_memory[36783] = 3'b111;
        rom_memory[36784] = 3'b111;
        rom_memory[36785] = 3'b110;
        rom_memory[36786] = 3'b000;
        rom_memory[36787] = 3'b000;
        rom_memory[36788] = 3'b000;
        rom_memory[36789] = 3'b111;
        rom_memory[36790] = 3'b111;
        rom_memory[36791] = 3'b111;
        rom_memory[36792] = 3'b111;
        rom_memory[36793] = 3'b111;
        rom_memory[36794] = 3'b111;
        rom_memory[36795] = 3'b111;
        rom_memory[36796] = 3'b111;
        rom_memory[36797] = 3'b110;
        rom_memory[36798] = 3'b110;
        rom_memory[36799] = 3'b110;
        rom_memory[36800] = 3'b111;
        rom_memory[36801] = 3'b000;
        rom_memory[36802] = 3'b000;
        rom_memory[36803] = 3'b000;
        rom_memory[36804] = 3'b000;
        rom_memory[36805] = 3'b000;
        rom_memory[36806] = 3'b000;
        rom_memory[36807] = 3'b000;
        rom_memory[36808] = 3'b000;
        rom_memory[36809] = 3'b111;
        rom_memory[36810] = 3'b000;
        rom_memory[36811] = 3'b111;
        rom_memory[36812] = 3'b111;
        rom_memory[36813] = 3'b000;
        rom_memory[36814] = 3'b000;
        rom_memory[36815] = 3'b000;
        rom_memory[36816] = 3'b110;
        rom_memory[36817] = 3'b110;
        rom_memory[36818] = 3'b110;
        rom_memory[36819] = 3'b110;
        rom_memory[36820] = 3'b110;
        rom_memory[36821] = 3'b110;
        rom_memory[36822] = 3'b110;
        rom_memory[36823] = 3'b110;
        rom_memory[36824] = 3'b110;
        rom_memory[36825] = 3'b110;
        rom_memory[36826] = 3'b110;
        rom_memory[36827] = 3'b110;
        rom_memory[36828] = 3'b110;
        rom_memory[36829] = 3'b110;
        rom_memory[36830] = 3'b110;
        rom_memory[36831] = 3'b110;
        rom_memory[36832] = 3'b110;
        rom_memory[36833] = 3'b110;
        rom_memory[36834] = 3'b110;
        rom_memory[36835] = 3'b110;
        rom_memory[36836] = 3'b110;
        rom_memory[36837] = 3'b110;
        rom_memory[36838] = 3'b110;
        rom_memory[36839] = 3'b110;
        rom_memory[36840] = 3'b110;
        rom_memory[36841] = 3'b110;
        rom_memory[36842] = 3'b110;
        rom_memory[36843] = 3'b110;
        rom_memory[36844] = 3'b110;
        rom_memory[36845] = 3'b110;
        rom_memory[36846] = 3'b110;
        rom_memory[36847] = 3'b110;
        rom_memory[36848] = 3'b110;
        rom_memory[36849] = 3'b110;
        rom_memory[36850] = 3'b110;
        rom_memory[36851] = 3'b110;
        rom_memory[36852] = 3'b110;
        rom_memory[36853] = 3'b110;
        rom_memory[36854] = 3'b110;
        rom_memory[36855] = 3'b110;
        rom_memory[36856] = 3'b110;
        rom_memory[36857] = 3'b110;
        rom_memory[36858] = 3'b110;
        rom_memory[36859] = 3'b110;
        rom_memory[36860] = 3'b110;
        rom_memory[36861] = 3'b110;
        rom_memory[36862] = 3'b110;
        rom_memory[36863] = 3'b110;
        rom_memory[36864] = 3'b110;
        rom_memory[36865] = 3'b110;
        rom_memory[36866] = 3'b110;
        rom_memory[36867] = 3'b110;
        rom_memory[36868] = 3'b110;
        rom_memory[36869] = 3'b110;
        rom_memory[36870] = 3'b110;
        rom_memory[36871] = 3'b110;
        rom_memory[36872] = 3'b110;
        rom_memory[36873] = 3'b000;
        rom_memory[36874] = 3'b000;
        rom_memory[36875] = 3'b000;
        rom_memory[36876] = 3'b000;
        rom_memory[36877] = 3'b000;
        rom_memory[36878] = 3'b110;
        rom_memory[36879] = 3'b111;
        rom_memory[36880] = 3'b000;
        rom_memory[36881] = 3'b000;
        rom_memory[36882] = 3'b100;
        rom_memory[36883] = 3'b000;
        rom_memory[36884] = 3'b000;
        rom_memory[36885] = 3'b000;
        rom_memory[36886] = 3'b000;
        rom_memory[36887] = 3'b100;
        rom_memory[36888] = 3'b111;
        rom_memory[36889] = 3'b110;
        rom_memory[36890] = 3'b110;
        rom_memory[36891] = 3'b110;
        rom_memory[36892] = 3'b110;
        rom_memory[36893] = 3'b110;
        rom_memory[36894] = 3'b110;
        rom_memory[36895] = 3'b110;
        rom_memory[36896] = 3'b110;
        rom_memory[36897] = 3'b110;
        rom_memory[36898] = 3'b110;
        rom_memory[36899] = 3'b110;
        rom_memory[36900] = 3'b110;
        rom_memory[36901] = 3'b110;
        rom_memory[36902] = 3'b110;
        rom_memory[36903] = 3'b110;
        rom_memory[36904] = 3'b110;
        rom_memory[36905] = 3'b110;
        rom_memory[36906] = 3'b110;
        rom_memory[36907] = 3'b110;
        rom_memory[36908] = 3'b110;
        rom_memory[36909] = 3'b110;
        rom_memory[36910] = 3'b110;
        rom_memory[36911] = 3'b110;
        rom_memory[36912] = 3'b110;
        rom_memory[36913] = 3'b110;
        rom_memory[36914] = 3'b110;
        rom_memory[36915] = 3'b110;
        rom_memory[36916] = 3'b110;
        rom_memory[36917] = 3'b110;
        rom_memory[36918] = 3'b110;
        rom_memory[36919] = 3'b111;
        rom_memory[36920] = 3'b111;
        rom_memory[36921] = 3'b111;
        rom_memory[36922] = 3'b111;
        rom_memory[36923] = 3'b111;
        rom_memory[36924] = 3'b111;
        rom_memory[36925] = 3'b111;
        rom_memory[36926] = 3'b111;
        rom_memory[36927] = 3'b111;
        rom_memory[36928] = 3'b111;
        rom_memory[36929] = 3'b111;
        rom_memory[36930] = 3'b111;
        rom_memory[36931] = 3'b111;
        rom_memory[36932] = 3'b111;
        rom_memory[36933] = 3'b111;
        rom_memory[36934] = 3'b111;
        rom_memory[36935] = 3'b111;
        rom_memory[36936] = 3'b111;
        rom_memory[36937] = 3'b111;
        rom_memory[36938] = 3'b111;
        rom_memory[36939] = 3'b111;
        rom_memory[36940] = 3'b111;
        rom_memory[36941] = 3'b111;
        rom_memory[36942] = 3'b111;
        rom_memory[36943] = 3'b111;
        rom_memory[36944] = 3'b111;
        rom_memory[36945] = 3'b111;
        rom_memory[36946] = 3'b111;
        rom_memory[36947] = 3'b111;
        rom_memory[36948] = 3'b111;
        rom_memory[36949] = 3'b111;
        rom_memory[36950] = 3'b111;
        rom_memory[36951] = 3'b111;
        rom_memory[36952] = 3'b111;
        rom_memory[36953] = 3'b111;
        rom_memory[36954] = 3'b111;
        rom_memory[36955] = 3'b111;
        rom_memory[36956] = 3'b111;
        rom_memory[36957] = 3'b111;
        rom_memory[36958] = 3'b111;
        rom_memory[36959] = 3'b111;
        rom_memory[36960] = 3'b110;
        rom_memory[36961] = 3'b110;
        rom_memory[36962] = 3'b110;
        rom_memory[36963] = 3'b110;
        rom_memory[36964] = 3'b110;
        rom_memory[36965] = 3'b110;
        rom_memory[36966] = 3'b110;
        rom_memory[36967] = 3'b111;
        rom_memory[36968] = 3'b111;
        rom_memory[36969] = 3'b111;
        rom_memory[36970] = 3'b111;
        rom_memory[36971] = 3'b111;
        rom_memory[36972] = 3'b111;
        rom_memory[36973] = 3'b111;
        rom_memory[36974] = 3'b111;
        rom_memory[36975] = 3'b111;
        rom_memory[36976] = 3'b111;
        rom_memory[36977] = 3'b111;
        rom_memory[36978] = 3'b111;
        rom_memory[36979] = 3'b111;
        rom_memory[36980] = 3'b111;
        rom_memory[36981] = 3'b111;
        rom_memory[36982] = 3'b111;
        rom_memory[36983] = 3'b111;
        rom_memory[36984] = 3'b110;
        rom_memory[36985] = 3'b110;
        rom_memory[36986] = 3'b110;
        rom_memory[36987] = 3'b110;
        rom_memory[36988] = 3'b110;
        rom_memory[36989] = 3'b110;
        rom_memory[36990] = 3'b110;
        rom_memory[36991] = 3'b110;
        rom_memory[36992] = 3'b110;
        rom_memory[36993] = 3'b110;
        rom_memory[36994] = 3'b110;
        rom_memory[36995] = 3'b110;
        rom_memory[36996] = 3'b110;
        rom_memory[36997] = 3'b110;
        rom_memory[36998] = 3'b110;
        rom_memory[36999] = 3'b110;
        rom_memory[37000] = 3'b110;
        rom_memory[37001] = 3'b110;
        rom_memory[37002] = 3'b111;
        rom_memory[37003] = 3'b111;
        rom_memory[37004] = 3'b111;
        rom_memory[37005] = 3'b111;
        rom_memory[37006] = 3'b111;
        rom_memory[37007] = 3'b111;
        rom_memory[37008] = 3'b111;
        rom_memory[37009] = 3'b111;
        rom_memory[37010] = 3'b111;
        rom_memory[37011] = 3'b110;
        rom_memory[37012] = 3'b110;
        rom_memory[37013] = 3'b110;
        rom_memory[37014] = 3'b110;
        rom_memory[37015] = 3'b010;
        rom_memory[37016] = 3'b000;
        rom_memory[37017] = 3'b110;
        rom_memory[37018] = 3'b110;
        rom_memory[37019] = 3'b110;
        rom_memory[37020] = 3'b110;
        rom_memory[37021] = 3'b110;
        rom_memory[37022] = 3'b111;
        rom_memory[37023] = 3'b111;
        rom_memory[37024] = 3'b111;
        rom_memory[37025] = 3'b110;
        rom_memory[37026] = 3'b000;
        rom_memory[37027] = 3'b000;
        rom_memory[37028] = 3'b000;
        rom_memory[37029] = 3'b111;
        rom_memory[37030] = 3'b100;
        rom_memory[37031] = 3'b111;
        rom_memory[37032] = 3'b111;
        rom_memory[37033] = 3'b111;
        rom_memory[37034] = 3'b110;
        rom_memory[37035] = 3'b111;
        rom_memory[37036] = 3'b111;
        rom_memory[37037] = 3'b111;
        rom_memory[37038] = 3'b110;
        rom_memory[37039] = 3'b110;
        rom_memory[37040] = 3'b110;
        rom_memory[37041] = 3'b000;
        rom_memory[37042] = 3'b000;
        rom_memory[37043] = 3'b000;
        rom_memory[37044] = 3'b000;
        rom_memory[37045] = 3'b000;
        rom_memory[37046] = 3'b000;
        rom_memory[37047] = 3'b000;
        rom_memory[37048] = 3'b111;
        rom_memory[37049] = 3'b111;
        rom_memory[37050] = 3'b111;
        rom_memory[37051] = 3'b111;
        rom_memory[37052] = 3'b111;
        rom_memory[37053] = 3'b111;
        rom_memory[37054] = 3'b000;
        rom_memory[37055] = 3'b000;
        rom_memory[37056] = 3'b110;
        rom_memory[37057] = 3'b110;
        rom_memory[37058] = 3'b110;
        rom_memory[37059] = 3'b110;
        rom_memory[37060] = 3'b110;
        rom_memory[37061] = 3'b110;
        rom_memory[37062] = 3'b110;
        rom_memory[37063] = 3'b110;
        rom_memory[37064] = 3'b110;
        rom_memory[37065] = 3'b110;
        rom_memory[37066] = 3'b110;
        rom_memory[37067] = 3'b110;
        rom_memory[37068] = 3'b110;
        rom_memory[37069] = 3'b110;
        rom_memory[37070] = 3'b110;
        rom_memory[37071] = 3'b110;
        rom_memory[37072] = 3'b110;
        rom_memory[37073] = 3'b110;
        rom_memory[37074] = 3'b110;
        rom_memory[37075] = 3'b110;
        rom_memory[37076] = 3'b110;
        rom_memory[37077] = 3'b110;
        rom_memory[37078] = 3'b110;
        rom_memory[37079] = 3'b110;
        rom_memory[37080] = 3'b110;
        rom_memory[37081] = 3'b110;
        rom_memory[37082] = 3'b110;
        rom_memory[37083] = 3'b110;
        rom_memory[37084] = 3'b110;
        rom_memory[37085] = 3'b110;
        rom_memory[37086] = 3'b110;
        rom_memory[37087] = 3'b110;
        rom_memory[37088] = 3'b110;
        rom_memory[37089] = 3'b110;
        rom_memory[37090] = 3'b110;
        rom_memory[37091] = 3'b110;
        rom_memory[37092] = 3'b110;
        rom_memory[37093] = 3'b110;
        rom_memory[37094] = 3'b110;
        rom_memory[37095] = 3'b110;
        rom_memory[37096] = 3'b110;
        rom_memory[37097] = 3'b110;
        rom_memory[37098] = 3'b110;
        rom_memory[37099] = 3'b110;
        rom_memory[37100] = 3'b110;
        rom_memory[37101] = 3'b110;
        rom_memory[37102] = 3'b110;
        rom_memory[37103] = 3'b110;
        rom_memory[37104] = 3'b110;
        rom_memory[37105] = 3'b110;
        rom_memory[37106] = 3'b110;
        rom_memory[37107] = 3'b110;
        rom_memory[37108] = 3'b110;
        rom_memory[37109] = 3'b110;
        rom_memory[37110] = 3'b110;
        rom_memory[37111] = 3'b110;
        rom_memory[37112] = 3'b110;
        rom_memory[37113] = 3'b110;
        rom_memory[37114] = 3'b000;
        rom_memory[37115] = 3'b000;
        rom_memory[37116] = 3'b000;
        rom_memory[37117] = 3'b000;
        rom_memory[37118] = 3'b000;
        rom_memory[37119] = 3'b110;
        rom_memory[37120] = 3'b111;
        rom_memory[37121] = 3'b000;
        rom_memory[37122] = 3'b000;
        rom_memory[37123] = 3'b100;
        rom_memory[37124] = 3'b000;
        rom_memory[37125] = 3'b000;
        rom_memory[37126] = 3'b000;
        rom_memory[37127] = 3'b000;
        rom_memory[37128] = 3'b000;
        rom_memory[37129] = 3'b111;
        rom_memory[37130] = 3'b111;
        rom_memory[37131] = 3'b110;
        rom_memory[37132] = 3'b110;
        rom_memory[37133] = 3'b110;
        rom_memory[37134] = 3'b110;
        rom_memory[37135] = 3'b110;
        rom_memory[37136] = 3'b110;
        rom_memory[37137] = 3'b110;
        rom_memory[37138] = 3'b110;
        rom_memory[37139] = 3'b110;
        rom_memory[37140] = 3'b110;
        rom_memory[37141] = 3'b110;
        rom_memory[37142] = 3'b110;
        rom_memory[37143] = 3'b110;
        rom_memory[37144] = 3'b110;
        rom_memory[37145] = 3'b110;
        rom_memory[37146] = 3'b110;
        rom_memory[37147] = 3'b110;
        rom_memory[37148] = 3'b110;
        rom_memory[37149] = 3'b110;
        rom_memory[37150] = 3'b110;
        rom_memory[37151] = 3'b110;
        rom_memory[37152] = 3'b110;
        rom_memory[37153] = 3'b110;
        rom_memory[37154] = 3'b110;
        rom_memory[37155] = 3'b110;
        rom_memory[37156] = 3'b110;
        rom_memory[37157] = 3'b110;
        rom_memory[37158] = 3'b110;
        rom_memory[37159] = 3'b110;
        rom_memory[37160] = 3'b111;
        rom_memory[37161] = 3'b111;
        rom_memory[37162] = 3'b111;
        rom_memory[37163] = 3'b111;
        rom_memory[37164] = 3'b111;
        rom_memory[37165] = 3'b111;
        rom_memory[37166] = 3'b111;
        rom_memory[37167] = 3'b111;
        rom_memory[37168] = 3'b111;
        rom_memory[37169] = 3'b111;
        rom_memory[37170] = 3'b111;
        rom_memory[37171] = 3'b111;
        rom_memory[37172] = 3'b111;
        rom_memory[37173] = 3'b111;
        rom_memory[37174] = 3'b111;
        rom_memory[37175] = 3'b111;
        rom_memory[37176] = 3'b111;
        rom_memory[37177] = 3'b111;
        rom_memory[37178] = 3'b111;
        rom_memory[37179] = 3'b111;
        rom_memory[37180] = 3'b111;
        rom_memory[37181] = 3'b111;
        rom_memory[37182] = 3'b111;
        rom_memory[37183] = 3'b111;
        rom_memory[37184] = 3'b111;
        rom_memory[37185] = 3'b111;
        rom_memory[37186] = 3'b111;
        rom_memory[37187] = 3'b111;
        rom_memory[37188] = 3'b111;
        rom_memory[37189] = 3'b111;
        rom_memory[37190] = 3'b111;
        rom_memory[37191] = 3'b111;
        rom_memory[37192] = 3'b111;
        rom_memory[37193] = 3'b111;
        rom_memory[37194] = 3'b111;
        rom_memory[37195] = 3'b111;
        rom_memory[37196] = 3'b111;
        rom_memory[37197] = 3'b111;
        rom_memory[37198] = 3'b111;
        rom_memory[37199] = 3'b111;
        rom_memory[37200] = 3'b110;
        rom_memory[37201] = 3'b110;
        rom_memory[37202] = 3'b110;
        rom_memory[37203] = 3'b110;
        rom_memory[37204] = 3'b110;
        rom_memory[37205] = 3'b110;
        rom_memory[37206] = 3'b110;
        rom_memory[37207] = 3'b111;
        rom_memory[37208] = 3'b111;
        rom_memory[37209] = 3'b111;
        rom_memory[37210] = 3'b111;
        rom_memory[37211] = 3'b111;
        rom_memory[37212] = 3'b111;
        rom_memory[37213] = 3'b111;
        rom_memory[37214] = 3'b111;
        rom_memory[37215] = 3'b111;
        rom_memory[37216] = 3'b111;
        rom_memory[37217] = 3'b111;
        rom_memory[37218] = 3'b111;
        rom_memory[37219] = 3'b111;
        rom_memory[37220] = 3'b111;
        rom_memory[37221] = 3'b111;
        rom_memory[37222] = 3'b111;
        rom_memory[37223] = 3'b111;
        rom_memory[37224] = 3'b110;
        rom_memory[37225] = 3'b110;
        rom_memory[37226] = 3'b110;
        rom_memory[37227] = 3'b110;
        rom_memory[37228] = 3'b110;
        rom_memory[37229] = 3'b110;
        rom_memory[37230] = 3'b110;
        rom_memory[37231] = 3'b110;
        rom_memory[37232] = 3'b110;
        rom_memory[37233] = 3'b110;
        rom_memory[37234] = 3'b110;
        rom_memory[37235] = 3'b110;
        rom_memory[37236] = 3'b110;
        rom_memory[37237] = 3'b110;
        rom_memory[37238] = 3'b110;
        rom_memory[37239] = 3'b110;
        rom_memory[37240] = 3'b110;
        rom_memory[37241] = 3'b110;
        rom_memory[37242] = 3'b110;
        rom_memory[37243] = 3'b111;
        rom_memory[37244] = 3'b111;
        rom_memory[37245] = 3'b111;
        rom_memory[37246] = 3'b111;
        rom_memory[37247] = 3'b111;
        rom_memory[37248] = 3'b111;
        rom_memory[37249] = 3'b111;
        rom_memory[37250] = 3'b111;
        rom_memory[37251] = 3'b111;
        rom_memory[37252] = 3'b111;
        rom_memory[37253] = 3'b110;
        rom_memory[37254] = 3'b110;
        rom_memory[37255] = 3'b110;
        rom_memory[37256] = 3'b000;
        rom_memory[37257] = 3'b000;
        rom_memory[37258] = 3'b000;
        rom_memory[37259] = 3'b110;
        rom_memory[37260] = 3'b110;
        rom_memory[37261] = 3'b110;
        rom_memory[37262] = 3'b111;
        rom_memory[37263] = 3'b111;
        rom_memory[37264] = 3'b111;
        rom_memory[37265] = 3'b110;
        rom_memory[37266] = 3'b000;
        rom_memory[37267] = 3'b000;
        rom_memory[37268] = 3'b000;
        rom_memory[37269] = 3'b111;
        rom_memory[37270] = 3'b000;
        rom_memory[37271] = 3'b110;
        rom_memory[37272] = 3'b111;
        rom_memory[37273] = 3'b111;
        rom_memory[37274] = 3'b111;
        rom_memory[37275] = 3'b110;
        rom_memory[37276] = 3'b111;
        rom_memory[37277] = 3'b111;
        rom_memory[37278] = 3'b111;
        rom_memory[37279] = 3'b110;
        rom_memory[37280] = 3'b110;
        rom_memory[37281] = 3'b000;
        rom_memory[37282] = 3'b000;
        rom_memory[37283] = 3'b000;
        rom_memory[37284] = 3'b000;
        rom_memory[37285] = 3'b001;
        rom_memory[37286] = 3'b011;
        rom_memory[37287] = 3'b111;
        rom_memory[37288] = 3'b111;
        rom_memory[37289] = 3'b111;
        rom_memory[37290] = 3'b111;
        rom_memory[37291] = 3'b111;
        rom_memory[37292] = 3'b111;
        rom_memory[37293] = 3'b111;
        rom_memory[37294] = 3'b001;
        rom_memory[37295] = 3'b000;
        rom_memory[37296] = 3'b111;
        rom_memory[37297] = 3'b111;
        rom_memory[37298] = 3'b110;
        rom_memory[37299] = 3'b110;
        rom_memory[37300] = 3'b110;
        rom_memory[37301] = 3'b110;
        rom_memory[37302] = 3'b110;
        rom_memory[37303] = 3'b110;
        rom_memory[37304] = 3'b110;
        rom_memory[37305] = 3'b110;
        rom_memory[37306] = 3'b110;
        rom_memory[37307] = 3'b110;
        rom_memory[37308] = 3'b110;
        rom_memory[37309] = 3'b110;
        rom_memory[37310] = 3'b110;
        rom_memory[37311] = 3'b110;
        rom_memory[37312] = 3'b110;
        rom_memory[37313] = 3'b110;
        rom_memory[37314] = 3'b110;
        rom_memory[37315] = 3'b110;
        rom_memory[37316] = 3'b110;
        rom_memory[37317] = 3'b110;
        rom_memory[37318] = 3'b110;
        rom_memory[37319] = 3'b110;
        rom_memory[37320] = 3'b110;
        rom_memory[37321] = 3'b110;
        rom_memory[37322] = 3'b110;
        rom_memory[37323] = 3'b110;
        rom_memory[37324] = 3'b110;
        rom_memory[37325] = 3'b110;
        rom_memory[37326] = 3'b110;
        rom_memory[37327] = 3'b110;
        rom_memory[37328] = 3'b110;
        rom_memory[37329] = 3'b110;
        rom_memory[37330] = 3'b110;
        rom_memory[37331] = 3'b110;
        rom_memory[37332] = 3'b110;
        rom_memory[37333] = 3'b110;
        rom_memory[37334] = 3'b110;
        rom_memory[37335] = 3'b110;
        rom_memory[37336] = 3'b110;
        rom_memory[37337] = 3'b110;
        rom_memory[37338] = 3'b110;
        rom_memory[37339] = 3'b110;
        rom_memory[37340] = 3'b110;
        rom_memory[37341] = 3'b110;
        rom_memory[37342] = 3'b110;
        rom_memory[37343] = 3'b110;
        rom_memory[37344] = 3'b110;
        rom_memory[37345] = 3'b110;
        rom_memory[37346] = 3'b110;
        rom_memory[37347] = 3'b110;
        rom_memory[37348] = 3'b110;
        rom_memory[37349] = 3'b110;
        rom_memory[37350] = 3'b110;
        rom_memory[37351] = 3'b110;
        rom_memory[37352] = 3'b110;
        rom_memory[37353] = 3'b110;
        rom_memory[37354] = 3'b110;
        rom_memory[37355] = 3'b000;
        rom_memory[37356] = 3'b000;
        rom_memory[37357] = 3'b000;
        rom_memory[37358] = 3'b000;
        rom_memory[37359] = 3'b000;
        rom_memory[37360] = 3'b110;
        rom_memory[37361] = 3'b111;
        rom_memory[37362] = 3'b000;
        rom_memory[37363] = 3'b000;
        rom_memory[37364] = 3'b100;
        rom_memory[37365] = 3'b000;
        rom_memory[37366] = 3'b000;
        rom_memory[37367] = 3'b000;
        rom_memory[37368] = 3'b000;
        rom_memory[37369] = 3'b000;
        rom_memory[37370] = 3'b110;
        rom_memory[37371] = 3'b111;
        rom_memory[37372] = 3'b110;
        rom_memory[37373] = 3'b110;
        rom_memory[37374] = 3'b110;
        rom_memory[37375] = 3'b110;
        rom_memory[37376] = 3'b110;
        rom_memory[37377] = 3'b110;
        rom_memory[37378] = 3'b110;
        rom_memory[37379] = 3'b110;
        rom_memory[37380] = 3'b110;
        rom_memory[37381] = 3'b110;
        rom_memory[37382] = 3'b110;
        rom_memory[37383] = 3'b110;
        rom_memory[37384] = 3'b110;
        rom_memory[37385] = 3'b110;
        rom_memory[37386] = 3'b110;
        rom_memory[37387] = 3'b110;
        rom_memory[37388] = 3'b110;
        rom_memory[37389] = 3'b110;
        rom_memory[37390] = 3'b110;
        rom_memory[37391] = 3'b110;
        rom_memory[37392] = 3'b110;
        rom_memory[37393] = 3'b110;
        rom_memory[37394] = 3'b110;
        rom_memory[37395] = 3'b110;
        rom_memory[37396] = 3'b110;
        rom_memory[37397] = 3'b110;
        rom_memory[37398] = 3'b110;
        rom_memory[37399] = 3'b110;
        rom_memory[37400] = 3'b110;
        rom_memory[37401] = 3'b111;
        rom_memory[37402] = 3'b111;
        rom_memory[37403] = 3'b111;
        rom_memory[37404] = 3'b111;
        rom_memory[37405] = 3'b111;
        rom_memory[37406] = 3'b111;
        rom_memory[37407] = 3'b111;
        rom_memory[37408] = 3'b111;
        rom_memory[37409] = 3'b111;
        rom_memory[37410] = 3'b111;
        rom_memory[37411] = 3'b111;
        rom_memory[37412] = 3'b111;
        rom_memory[37413] = 3'b111;
        rom_memory[37414] = 3'b111;
        rom_memory[37415] = 3'b111;
        rom_memory[37416] = 3'b111;
        rom_memory[37417] = 3'b111;
        rom_memory[37418] = 3'b111;
        rom_memory[37419] = 3'b111;
        rom_memory[37420] = 3'b111;
        rom_memory[37421] = 3'b111;
        rom_memory[37422] = 3'b111;
        rom_memory[37423] = 3'b111;
        rom_memory[37424] = 3'b111;
        rom_memory[37425] = 3'b111;
        rom_memory[37426] = 3'b111;
        rom_memory[37427] = 3'b111;
        rom_memory[37428] = 3'b111;
        rom_memory[37429] = 3'b111;
        rom_memory[37430] = 3'b111;
        rom_memory[37431] = 3'b111;
        rom_memory[37432] = 3'b111;
        rom_memory[37433] = 3'b111;
        rom_memory[37434] = 3'b111;
        rom_memory[37435] = 3'b111;
        rom_memory[37436] = 3'b111;
        rom_memory[37437] = 3'b111;
        rom_memory[37438] = 3'b111;
        rom_memory[37439] = 3'b111;
        rom_memory[37440] = 3'b110;
        rom_memory[37441] = 3'b110;
        rom_memory[37442] = 3'b110;
        rom_memory[37443] = 3'b110;
        rom_memory[37444] = 3'b110;
        rom_memory[37445] = 3'b110;
        rom_memory[37446] = 3'b110;
        rom_memory[37447] = 3'b110;
        rom_memory[37448] = 3'b111;
        rom_memory[37449] = 3'b111;
        rom_memory[37450] = 3'b111;
        rom_memory[37451] = 3'b111;
        rom_memory[37452] = 3'b111;
        rom_memory[37453] = 3'b111;
        rom_memory[37454] = 3'b111;
        rom_memory[37455] = 3'b111;
        rom_memory[37456] = 3'b111;
        rom_memory[37457] = 3'b111;
        rom_memory[37458] = 3'b111;
        rom_memory[37459] = 3'b111;
        rom_memory[37460] = 3'b111;
        rom_memory[37461] = 3'b111;
        rom_memory[37462] = 3'b111;
        rom_memory[37463] = 3'b111;
        rom_memory[37464] = 3'b110;
        rom_memory[37465] = 3'b110;
        rom_memory[37466] = 3'b110;
        rom_memory[37467] = 3'b110;
        rom_memory[37468] = 3'b110;
        rom_memory[37469] = 3'b110;
        rom_memory[37470] = 3'b110;
        rom_memory[37471] = 3'b110;
        rom_memory[37472] = 3'b110;
        rom_memory[37473] = 3'b110;
        rom_memory[37474] = 3'b110;
        rom_memory[37475] = 3'b110;
        rom_memory[37476] = 3'b110;
        rom_memory[37477] = 3'b110;
        rom_memory[37478] = 3'b110;
        rom_memory[37479] = 3'b110;
        rom_memory[37480] = 3'b110;
        rom_memory[37481] = 3'b110;
        rom_memory[37482] = 3'b110;
        rom_memory[37483] = 3'b111;
        rom_memory[37484] = 3'b111;
        rom_memory[37485] = 3'b111;
        rom_memory[37486] = 3'b111;
        rom_memory[37487] = 3'b111;
        rom_memory[37488] = 3'b111;
        rom_memory[37489] = 3'b111;
        rom_memory[37490] = 3'b111;
        rom_memory[37491] = 3'b111;
        rom_memory[37492] = 3'b111;
        rom_memory[37493] = 3'b111;
        rom_memory[37494] = 3'b111;
        rom_memory[37495] = 3'b110;
        rom_memory[37496] = 3'b000;
        rom_memory[37497] = 3'b000;
        rom_memory[37498] = 3'b000;
        rom_memory[37499] = 3'b110;
        rom_memory[37500] = 3'b110;
        rom_memory[37501] = 3'b110;
        rom_memory[37502] = 3'b111;
        rom_memory[37503] = 3'b111;
        rom_memory[37504] = 3'b110;
        rom_memory[37505] = 3'b111;
        rom_memory[37506] = 3'b000;
        rom_memory[37507] = 3'b000;
        rom_memory[37508] = 3'b000;
        rom_memory[37509] = 3'b000;
        rom_memory[37510] = 3'b000;
        rom_memory[37511] = 3'b110;
        rom_memory[37512] = 3'b110;
        rom_memory[37513] = 3'b110;
        rom_memory[37514] = 3'b111;
        rom_memory[37515] = 3'b110;
        rom_memory[37516] = 3'b111;
        rom_memory[37517] = 3'b111;
        rom_memory[37518] = 3'b111;
        rom_memory[37519] = 3'b111;
        rom_memory[37520] = 3'b110;
        rom_memory[37521] = 3'b000;
        rom_memory[37522] = 3'b000;
        rom_memory[37523] = 3'b000;
        rom_memory[37524] = 3'b011;
        rom_memory[37525] = 3'b011;
        rom_memory[37526] = 3'b111;
        rom_memory[37527] = 3'b111;
        rom_memory[37528] = 3'b111;
        rom_memory[37529] = 3'b111;
        rom_memory[37530] = 3'b111;
        rom_memory[37531] = 3'b111;
        rom_memory[37532] = 3'b111;
        rom_memory[37533] = 3'b111;
        rom_memory[37534] = 3'b001;
        rom_memory[37535] = 3'b001;
        rom_memory[37536] = 3'b011;
        rom_memory[37537] = 3'b111;
        rom_memory[37538] = 3'b111;
        rom_memory[37539] = 3'b111;
        rom_memory[37540] = 3'b110;
        rom_memory[37541] = 3'b110;
        rom_memory[37542] = 3'b110;
        rom_memory[37543] = 3'b110;
        rom_memory[37544] = 3'b110;
        rom_memory[37545] = 3'b110;
        rom_memory[37546] = 3'b110;
        rom_memory[37547] = 3'b110;
        rom_memory[37548] = 3'b110;
        rom_memory[37549] = 3'b110;
        rom_memory[37550] = 3'b110;
        rom_memory[37551] = 3'b110;
        rom_memory[37552] = 3'b110;
        rom_memory[37553] = 3'b110;
        rom_memory[37554] = 3'b110;
        rom_memory[37555] = 3'b110;
        rom_memory[37556] = 3'b110;
        rom_memory[37557] = 3'b110;
        rom_memory[37558] = 3'b110;
        rom_memory[37559] = 3'b110;
        rom_memory[37560] = 3'b110;
        rom_memory[37561] = 3'b110;
        rom_memory[37562] = 3'b110;
        rom_memory[37563] = 3'b110;
        rom_memory[37564] = 3'b110;
        rom_memory[37565] = 3'b110;
        rom_memory[37566] = 3'b110;
        rom_memory[37567] = 3'b110;
        rom_memory[37568] = 3'b110;
        rom_memory[37569] = 3'b110;
        rom_memory[37570] = 3'b110;
        rom_memory[37571] = 3'b110;
        rom_memory[37572] = 3'b110;
        rom_memory[37573] = 3'b110;
        rom_memory[37574] = 3'b110;
        rom_memory[37575] = 3'b110;
        rom_memory[37576] = 3'b110;
        rom_memory[37577] = 3'b110;
        rom_memory[37578] = 3'b110;
        rom_memory[37579] = 3'b110;
        rom_memory[37580] = 3'b110;
        rom_memory[37581] = 3'b110;
        rom_memory[37582] = 3'b110;
        rom_memory[37583] = 3'b110;
        rom_memory[37584] = 3'b110;
        rom_memory[37585] = 3'b110;
        rom_memory[37586] = 3'b110;
        rom_memory[37587] = 3'b110;
        rom_memory[37588] = 3'b110;
        rom_memory[37589] = 3'b110;
        rom_memory[37590] = 3'b110;
        rom_memory[37591] = 3'b110;
        rom_memory[37592] = 3'b110;
        rom_memory[37593] = 3'b110;
        rom_memory[37594] = 3'b110;
        rom_memory[37595] = 3'b111;
        rom_memory[37596] = 3'b110;
        rom_memory[37597] = 3'b000;
        rom_memory[37598] = 3'b000;
        rom_memory[37599] = 3'b000;
        rom_memory[37600] = 3'b000;
        rom_memory[37601] = 3'b110;
        rom_memory[37602] = 3'b111;
        rom_memory[37603] = 3'b000;
        rom_memory[37604] = 3'b000;
        rom_memory[37605] = 3'b000;
        rom_memory[37606] = 3'b000;
        rom_memory[37607] = 3'b000;
        rom_memory[37608] = 3'b000;
        rom_memory[37609] = 3'b000;
        rom_memory[37610] = 3'b000;
        rom_memory[37611] = 3'b110;
        rom_memory[37612] = 3'b111;
        rom_memory[37613] = 3'b110;
        rom_memory[37614] = 3'b110;
        rom_memory[37615] = 3'b110;
        rom_memory[37616] = 3'b110;
        rom_memory[37617] = 3'b110;
        rom_memory[37618] = 3'b110;
        rom_memory[37619] = 3'b110;
        rom_memory[37620] = 3'b110;
        rom_memory[37621] = 3'b110;
        rom_memory[37622] = 3'b110;
        rom_memory[37623] = 3'b110;
        rom_memory[37624] = 3'b110;
        rom_memory[37625] = 3'b110;
        rom_memory[37626] = 3'b110;
        rom_memory[37627] = 3'b110;
        rom_memory[37628] = 3'b110;
        rom_memory[37629] = 3'b110;
        rom_memory[37630] = 3'b110;
        rom_memory[37631] = 3'b110;
        rom_memory[37632] = 3'b110;
        rom_memory[37633] = 3'b110;
        rom_memory[37634] = 3'b110;
        rom_memory[37635] = 3'b110;
        rom_memory[37636] = 3'b110;
        rom_memory[37637] = 3'b110;
        rom_memory[37638] = 3'b110;
        rom_memory[37639] = 3'b110;
        rom_memory[37640] = 3'b110;
        rom_memory[37641] = 3'b111;
        rom_memory[37642] = 3'b111;
        rom_memory[37643] = 3'b111;
        rom_memory[37644] = 3'b111;
        rom_memory[37645] = 3'b111;
        rom_memory[37646] = 3'b111;
        rom_memory[37647] = 3'b111;
        rom_memory[37648] = 3'b111;
        rom_memory[37649] = 3'b111;
        rom_memory[37650] = 3'b111;
        rom_memory[37651] = 3'b111;
        rom_memory[37652] = 3'b111;
        rom_memory[37653] = 3'b111;
        rom_memory[37654] = 3'b111;
        rom_memory[37655] = 3'b111;
        rom_memory[37656] = 3'b111;
        rom_memory[37657] = 3'b111;
        rom_memory[37658] = 3'b111;
        rom_memory[37659] = 3'b111;
        rom_memory[37660] = 3'b111;
        rom_memory[37661] = 3'b111;
        rom_memory[37662] = 3'b111;
        rom_memory[37663] = 3'b111;
        rom_memory[37664] = 3'b111;
        rom_memory[37665] = 3'b111;
        rom_memory[37666] = 3'b111;
        rom_memory[37667] = 3'b111;
        rom_memory[37668] = 3'b111;
        rom_memory[37669] = 3'b111;
        rom_memory[37670] = 3'b111;
        rom_memory[37671] = 3'b111;
        rom_memory[37672] = 3'b111;
        rom_memory[37673] = 3'b111;
        rom_memory[37674] = 3'b111;
        rom_memory[37675] = 3'b111;
        rom_memory[37676] = 3'b111;
        rom_memory[37677] = 3'b111;
        rom_memory[37678] = 3'b111;
        rom_memory[37679] = 3'b111;
        rom_memory[37680] = 3'b110;
        rom_memory[37681] = 3'b110;
        rom_memory[37682] = 3'b110;
        rom_memory[37683] = 3'b110;
        rom_memory[37684] = 3'b110;
        rom_memory[37685] = 3'b110;
        rom_memory[37686] = 3'b110;
        rom_memory[37687] = 3'b110;
        rom_memory[37688] = 3'b111;
        rom_memory[37689] = 3'b111;
        rom_memory[37690] = 3'b111;
        rom_memory[37691] = 3'b111;
        rom_memory[37692] = 3'b111;
        rom_memory[37693] = 3'b111;
        rom_memory[37694] = 3'b111;
        rom_memory[37695] = 3'b111;
        rom_memory[37696] = 3'b111;
        rom_memory[37697] = 3'b111;
        rom_memory[37698] = 3'b111;
        rom_memory[37699] = 3'b111;
        rom_memory[37700] = 3'b111;
        rom_memory[37701] = 3'b111;
        rom_memory[37702] = 3'b111;
        rom_memory[37703] = 3'b111;
        rom_memory[37704] = 3'b111;
        rom_memory[37705] = 3'b110;
        rom_memory[37706] = 3'b110;
        rom_memory[37707] = 3'b110;
        rom_memory[37708] = 3'b110;
        rom_memory[37709] = 3'b110;
        rom_memory[37710] = 3'b110;
        rom_memory[37711] = 3'b110;
        rom_memory[37712] = 3'b110;
        rom_memory[37713] = 3'b110;
        rom_memory[37714] = 3'b110;
        rom_memory[37715] = 3'b110;
        rom_memory[37716] = 3'b110;
        rom_memory[37717] = 3'b110;
        rom_memory[37718] = 3'b110;
        rom_memory[37719] = 3'b110;
        rom_memory[37720] = 3'b110;
        rom_memory[37721] = 3'b110;
        rom_memory[37722] = 3'b110;
        rom_memory[37723] = 3'b111;
        rom_memory[37724] = 3'b111;
        rom_memory[37725] = 3'b111;
        rom_memory[37726] = 3'b111;
        rom_memory[37727] = 3'b111;
        rom_memory[37728] = 3'b111;
        rom_memory[37729] = 3'b111;
        rom_memory[37730] = 3'b111;
        rom_memory[37731] = 3'b111;
        rom_memory[37732] = 3'b111;
        rom_memory[37733] = 3'b111;
        rom_memory[37734] = 3'b111;
        rom_memory[37735] = 3'b111;
        rom_memory[37736] = 3'b111;
        rom_memory[37737] = 3'b110;
        rom_memory[37738] = 3'b110;
        rom_memory[37739] = 3'b110;
        rom_memory[37740] = 3'b110;
        rom_memory[37741] = 3'b110;
        rom_memory[37742] = 3'b111;
        rom_memory[37743] = 3'b111;
        rom_memory[37744] = 3'b110;
        rom_memory[37745] = 3'b000;
        rom_memory[37746] = 3'b110;
        rom_memory[37747] = 3'b100;
        rom_memory[37748] = 3'b000;
        rom_memory[37749] = 3'b000;
        rom_memory[37750] = 3'b000;
        rom_memory[37751] = 3'b110;
        rom_memory[37752] = 3'b110;
        rom_memory[37753] = 3'b110;
        rom_memory[37754] = 3'b111;
        rom_memory[37755] = 3'b110;
        rom_memory[37756] = 3'b110;
        rom_memory[37757] = 3'b110;
        rom_memory[37758] = 3'b111;
        rom_memory[37759] = 3'b111;
        rom_memory[37760] = 3'b000;
        rom_memory[37761] = 3'b000;
        rom_memory[37762] = 3'b000;
        rom_memory[37763] = 3'b000;
        rom_memory[37764] = 3'b111;
        rom_memory[37765] = 3'b100;
        rom_memory[37766] = 3'b100;
        rom_memory[37767] = 3'b111;
        rom_memory[37768] = 3'b110;
        rom_memory[37769] = 3'b110;
        rom_memory[37770] = 3'b111;
        rom_memory[37771] = 3'b111;
        rom_memory[37772] = 3'b111;
        rom_memory[37773] = 3'b111;
        rom_memory[37774] = 3'b001;
        rom_memory[37775] = 3'b001;
        rom_memory[37776] = 3'b011;
        rom_memory[37777] = 3'b111;
        rom_memory[37778] = 3'b111;
        rom_memory[37779] = 3'b111;
        rom_memory[37780] = 3'b111;
        rom_memory[37781] = 3'b110;
        rom_memory[37782] = 3'b110;
        rom_memory[37783] = 3'b110;
        rom_memory[37784] = 3'b110;
        rom_memory[37785] = 3'b110;
        rom_memory[37786] = 3'b110;
        rom_memory[37787] = 3'b110;
        rom_memory[37788] = 3'b110;
        rom_memory[37789] = 3'b110;
        rom_memory[37790] = 3'b110;
        rom_memory[37791] = 3'b110;
        rom_memory[37792] = 3'b110;
        rom_memory[37793] = 3'b110;
        rom_memory[37794] = 3'b110;
        rom_memory[37795] = 3'b110;
        rom_memory[37796] = 3'b110;
        rom_memory[37797] = 3'b110;
        rom_memory[37798] = 3'b110;
        rom_memory[37799] = 3'b110;
        rom_memory[37800] = 3'b110;
        rom_memory[37801] = 3'b110;
        rom_memory[37802] = 3'b110;
        rom_memory[37803] = 3'b110;
        rom_memory[37804] = 3'b110;
        rom_memory[37805] = 3'b110;
        rom_memory[37806] = 3'b110;
        rom_memory[37807] = 3'b110;
        rom_memory[37808] = 3'b110;
        rom_memory[37809] = 3'b110;
        rom_memory[37810] = 3'b110;
        rom_memory[37811] = 3'b110;
        rom_memory[37812] = 3'b110;
        rom_memory[37813] = 3'b110;
        rom_memory[37814] = 3'b110;
        rom_memory[37815] = 3'b110;
        rom_memory[37816] = 3'b110;
        rom_memory[37817] = 3'b110;
        rom_memory[37818] = 3'b110;
        rom_memory[37819] = 3'b110;
        rom_memory[37820] = 3'b110;
        rom_memory[37821] = 3'b110;
        rom_memory[37822] = 3'b110;
        rom_memory[37823] = 3'b110;
        rom_memory[37824] = 3'b110;
        rom_memory[37825] = 3'b110;
        rom_memory[37826] = 3'b110;
        rom_memory[37827] = 3'b110;
        rom_memory[37828] = 3'b110;
        rom_memory[37829] = 3'b110;
        rom_memory[37830] = 3'b110;
        rom_memory[37831] = 3'b110;
        rom_memory[37832] = 3'b110;
        rom_memory[37833] = 3'b110;
        rom_memory[37834] = 3'b110;
        rom_memory[37835] = 3'b110;
        rom_memory[37836] = 3'b111;
        rom_memory[37837] = 3'b110;
        rom_memory[37838] = 3'b000;
        rom_memory[37839] = 3'b000;
        rom_memory[37840] = 3'b000;
        rom_memory[37841] = 3'b000;
        rom_memory[37842] = 3'b110;
        rom_memory[37843] = 3'b111;
        rom_memory[37844] = 3'b000;
        rom_memory[37845] = 3'b000;
        rom_memory[37846] = 3'b000;
        rom_memory[37847] = 3'b000;
        rom_memory[37848] = 3'b000;
        rom_memory[37849] = 3'b000;
        rom_memory[37850] = 3'b000;
        rom_memory[37851] = 3'b000;
        rom_memory[37852] = 3'b110;
        rom_memory[37853] = 3'b111;
        rom_memory[37854] = 3'b110;
        rom_memory[37855] = 3'b110;
        rom_memory[37856] = 3'b110;
        rom_memory[37857] = 3'b110;
        rom_memory[37858] = 3'b110;
        rom_memory[37859] = 3'b110;
        rom_memory[37860] = 3'b110;
        rom_memory[37861] = 3'b110;
        rom_memory[37862] = 3'b110;
        rom_memory[37863] = 3'b110;
        rom_memory[37864] = 3'b110;
        rom_memory[37865] = 3'b110;
        rom_memory[37866] = 3'b110;
        rom_memory[37867] = 3'b110;
        rom_memory[37868] = 3'b110;
        rom_memory[37869] = 3'b110;
        rom_memory[37870] = 3'b110;
        rom_memory[37871] = 3'b110;
        rom_memory[37872] = 3'b110;
        rom_memory[37873] = 3'b110;
        rom_memory[37874] = 3'b110;
        rom_memory[37875] = 3'b110;
        rom_memory[37876] = 3'b110;
        rom_memory[37877] = 3'b110;
        rom_memory[37878] = 3'b110;
        rom_memory[37879] = 3'b110;
        rom_memory[37880] = 3'b110;
        rom_memory[37881] = 3'b110;
        rom_memory[37882] = 3'b110;
        rom_memory[37883] = 3'b110;
        rom_memory[37884] = 3'b111;
        rom_memory[37885] = 3'b111;
        rom_memory[37886] = 3'b111;
        rom_memory[37887] = 3'b111;
        rom_memory[37888] = 3'b111;
        rom_memory[37889] = 3'b111;
        rom_memory[37890] = 3'b111;
        rom_memory[37891] = 3'b111;
        rom_memory[37892] = 3'b111;
        rom_memory[37893] = 3'b111;
        rom_memory[37894] = 3'b111;
        rom_memory[37895] = 3'b111;
        rom_memory[37896] = 3'b111;
        rom_memory[37897] = 3'b111;
        rom_memory[37898] = 3'b111;
        rom_memory[37899] = 3'b111;
        rom_memory[37900] = 3'b111;
        rom_memory[37901] = 3'b111;
        rom_memory[37902] = 3'b111;
        rom_memory[37903] = 3'b111;
        rom_memory[37904] = 3'b111;
        rom_memory[37905] = 3'b111;
        rom_memory[37906] = 3'b111;
        rom_memory[37907] = 3'b111;
        rom_memory[37908] = 3'b111;
        rom_memory[37909] = 3'b111;
        rom_memory[37910] = 3'b111;
        rom_memory[37911] = 3'b111;
        rom_memory[37912] = 3'b111;
        rom_memory[37913] = 3'b111;
        rom_memory[37914] = 3'b111;
        rom_memory[37915] = 3'b111;
        rom_memory[37916] = 3'b111;
        rom_memory[37917] = 3'b111;
        rom_memory[37918] = 3'b111;
        rom_memory[37919] = 3'b111;
        rom_memory[37920] = 3'b110;
        rom_memory[37921] = 3'b110;
        rom_memory[37922] = 3'b110;
        rom_memory[37923] = 3'b110;
        rom_memory[37924] = 3'b110;
        rom_memory[37925] = 3'b110;
        rom_memory[37926] = 3'b110;
        rom_memory[37927] = 3'b110;
        rom_memory[37928] = 3'b110;
        rom_memory[37929] = 3'b111;
        rom_memory[37930] = 3'b111;
        rom_memory[37931] = 3'b111;
        rom_memory[37932] = 3'b111;
        rom_memory[37933] = 3'b111;
        rom_memory[37934] = 3'b111;
        rom_memory[37935] = 3'b111;
        rom_memory[37936] = 3'b111;
        rom_memory[37937] = 3'b111;
        rom_memory[37938] = 3'b111;
        rom_memory[37939] = 3'b111;
        rom_memory[37940] = 3'b111;
        rom_memory[37941] = 3'b111;
        rom_memory[37942] = 3'b111;
        rom_memory[37943] = 3'b111;
        rom_memory[37944] = 3'b111;
        rom_memory[37945] = 3'b110;
        rom_memory[37946] = 3'b110;
        rom_memory[37947] = 3'b110;
        rom_memory[37948] = 3'b110;
        rom_memory[37949] = 3'b110;
        rom_memory[37950] = 3'b110;
        rom_memory[37951] = 3'b110;
        rom_memory[37952] = 3'b110;
        rom_memory[37953] = 3'b110;
        rom_memory[37954] = 3'b110;
        rom_memory[37955] = 3'b110;
        rom_memory[37956] = 3'b110;
        rom_memory[37957] = 3'b110;
        rom_memory[37958] = 3'b110;
        rom_memory[37959] = 3'b110;
        rom_memory[37960] = 3'b110;
        rom_memory[37961] = 3'b110;
        rom_memory[37962] = 3'b110;
        rom_memory[37963] = 3'b111;
        rom_memory[37964] = 3'b111;
        rom_memory[37965] = 3'b111;
        rom_memory[37966] = 3'b111;
        rom_memory[37967] = 3'b111;
        rom_memory[37968] = 3'b111;
        rom_memory[37969] = 3'b111;
        rom_memory[37970] = 3'b111;
        rom_memory[37971] = 3'b111;
        rom_memory[37972] = 3'b111;
        rom_memory[37973] = 3'b111;
        rom_memory[37974] = 3'b111;
        rom_memory[37975] = 3'b111;
        rom_memory[37976] = 3'b111;
        rom_memory[37977] = 3'b111;
        rom_memory[37978] = 3'b111;
        rom_memory[37979] = 3'b111;
        rom_memory[37980] = 3'b110;
        rom_memory[37981] = 3'b110;
        rom_memory[37982] = 3'b111;
        rom_memory[37983] = 3'b111;
        rom_memory[37984] = 3'b110;
        rom_memory[37985] = 3'b100;
        rom_memory[37986] = 3'b110;
        rom_memory[37987] = 3'b000;
        rom_memory[37988] = 3'b000;
        rom_memory[37989] = 3'b000;
        rom_memory[37990] = 3'b000;
        rom_memory[37991] = 3'b110;
        rom_memory[37992] = 3'b110;
        rom_memory[37993] = 3'b110;
        rom_memory[37994] = 3'b110;
        rom_memory[37995] = 3'b111;
        rom_memory[37996] = 3'b110;
        rom_memory[37997] = 3'b110;
        rom_memory[37998] = 3'b111;
        rom_memory[37999] = 3'b111;
        rom_memory[38000] = 3'b111;
        rom_memory[38001] = 3'b000;
        rom_memory[38002] = 3'b000;
        rom_memory[38003] = 3'b111;
        rom_memory[38004] = 3'b111;
        rom_memory[38005] = 3'b100;
        rom_memory[38006] = 3'b110;
        rom_memory[38007] = 3'b100;
        rom_memory[38008] = 3'b100;
        rom_memory[38009] = 3'b110;
        rom_memory[38010] = 3'b111;
        rom_memory[38011] = 3'b111;
        rom_memory[38012] = 3'b111;
        rom_memory[38013] = 3'b111;
        rom_memory[38014] = 3'b011;
        rom_memory[38015] = 3'b011;
        rom_memory[38016] = 3'b011;
        rom_memory[38017] = 3'b111;
        rom_memory[38018] = 3'b111;
        rom_memory[38019] = 3'b111;
        rom_memory[38020] = 3'b111;
        rom_memory[38021] = 3'b110;
        rom_memory[38022] = 3'b110;
        rom_memory[38023] = 3'b110;
        rom_memory[38024] = 3'b110;
        rom_memory[38025] = 3'b110;
        rom_memory[38026] = 3'b110;
        rom_memory[38027] = 3'b110;
        rom_memory[38028] = 3'b110;
        rom_memory[38029] = 3'b110;
        rom_memory[38030] = 3'b110;
        rom_memory[38031] = 3'b110;
        rom_memory[38032] = 3'b110;
        rom_memory[38033] = 3'b110;
        rom_memory[38034] = 3'b110;
        rom_memory[38035] = 3'b110;
        rom_memory[38036] = 3'b110;
        rom_memory[38037] = 3'b110;
        rom_memory[38038] = 3'b110;
        rom_memory[38039] = 3'b110;
        rom_memory[38040] = 3'b110;
        rom_memory[38041] = 3'b110;
        rom_memory[38042] = 3'b110;
        rom_memory[38043] = 3'b110;
        rom_memory[38044] = 3'b110;
        rom_memory[38045] = 3'b110;
        rom_memory[38046] = 3'b110;
        rom_memory[38047] = 3'b110;
        rom_memory[38048] = 3'b110;
        rom_memory[38049] = 3'b110;
        rom_memory[38050] = 3'b110;
        rom_memory[38051] = 3'b110;
        rom_memory[38052] = 3'b110;
        rom_memory[38053] = 3'b110;
        rom_memory[38054] = 3'b110;
        rom_memory[38055] = 3'b110;
        rom_memory[38056] = 3'b110;
        rom_memory[38057] = 3'b110;
        rom_memory[38058] = 3'b110;
        rom_memory[38059] = 3'b110;
        rom_memory[38060] = 3'b110;
        rom_memory[38061] = 3'b110;
        rom_memory[38062] = 3'b110;
        rom_memory[38063] = 3'b110;
        rom_memory[38064] = 3'b110;
        rom_memory[38065] = 3'b110;
        rom_memory[38066] = 3'b110;
        rom_memory[38067] = 3'b110;
        rom_memory[38068] = 3'b110;
        rom_memory[38069] = 3'b110;
        rom_memory[38070] = 3'b110;
        rom_memory[38071] = 3'b110;
        rom_memory[38072] = 3'b110;
        rom_memory[38073] = 3'b110;
        rom_memory[38074] = 3'b110;
        rom_memory[38075] = 3'b110;
        rom_memory[38076] = 3'b110;
        rom_memory[38077] = 3'b111;
        rom_memory[38078] = 3'b110;
        rom_memory[38079] = 3'b000;
        rom_memory[38080] = 3'b000;
        rom_memory[38081] = 3'b000;
        rom_memory[38082] = 3'b000;
        rom_memory[38083] = 3'b100;
        rom_memory[38084] = 3'b110;
        rom_memory[38085] = 3'b000;
        rom_memory[38086] = 3'b000;
        rom_memory[38087] = 3'b000;
        rom_memory[38088] = 3'b000;
        rom_memory[38089] = 3'b000;
        rom_memory[38090] = 3'b000;
        rom_memory[38091] = 3'b000;
        rom_memory[38092] = 3'b000;
        rom_memory[38093] = 3'b110;
        rom_memory[38094] = 3'b111;
        rom_memory[38095] = 3'b110;
        rom_memory[38096] = 3'b110;
        rom_memory[38097] = 3'b110;
        rom_memory[38098] = 3'b110;
        rom_memory[38099] = 3'b110;
        rom_memory[38100] = 3'b110;
        rom_memory[38101] = 3'b110;
        rom_memory[38102] = 3'b110;
        rom_memory[38103] = 3'b110;
        rom_memory[38104] = 3'b110;
        rom_memory[38105] = 3'b110;
        rom_memory[38106] = 3'b110;
        rom_memory[38107] = 3'b110;
        rom_memory[38108] = 3'b110;
        rom_memory[38109] = 3'b110;
        rom_memory[38110] = 3'b110;
        rom_memory[38111] = 3'b110;
        rom_memory[38112] = 3'b110;
        rom_memory[38113] = 3'b110;
        rom_memory[38114] = 3'b110;
        rom_memory[38115] = 3'b110;
        rom_memory[38116] = 3'b110;
        rom_memory[38117] = 3'b110;
        rom_memory[38118] = 3'b110;
        rom_memory[38119] = 3'b110;
        rom_memory[38120] = 3'b110;
        rom_memory[38121] = 3'b110;
        rom_memory[38122] = 3'b110;
        rom_memory[38123] = 3'b110;
        rom_memory[38124] = 3'b111;
        rom_memory[38125] = 3'b111;
        rom_memory[38126] = 3'b111;
        rom_memory[38127] = 3'b111;
        rom_memory[38128] = 3'b111;
        rom_memory[38129] = 3'b111;
        rom_memory[38130] = 3'b111;
        rom_memory[38131] = 3'b111;
        rom_memory[38132] = 3'b111;
        rom_memory[38133] = 3'b111;
        rom_memory[38134] = 3'b111;
        rom_memory[38135] = 3'b111;
        rom_memory[38136] = 3'b111;
        rom_memory[38137] = 3'b111;
        rom_memory[38138] = 3'b111;
        rom_memory[38139] = 3'b111;
        rom_memory[38140] = 3'b111;
        rom_memory[38141] = 3'b111;
        rom_memory[38142] = 3'b111;
        rom_memory[38143] = 3'b111;
        rom_memory[38144] = 3'b111;
        rom_memory[38145] = 3'b111;
        rom_memory[38146] = 3'b111;
        rom_memory[38147] = 3'b111;
        rom_memory[38148] = 3'b111;
        rom_memory[38149] = 3'b111;
        rom_memory[38150] = 3'b111;
        rom_memory[38151] = 3'b111;
        rom_memory[38152] = 3'b111;
        rom_memory[38153] = 3'b111;
        rom_memory[38154] = 3'b111;
        rom_memory[38155] = 3'b111;
        rom_memory[38156] = 3'b111;
        rom_memory[38157] = 3'b111;
        rom_memory[38158] = 3'b111;
        rom_memory[38159] = 3'b111;
        rom_memory[38160] = 3'b110;
        rom_memory[38161] = 3'b110;
        rom_memory[38162] = 3'b110;
        rom_memory[38163] = 3'b110;
        rom_memory[38164] = 3'b110;
        rom_memory[38165] = 3'b110;
        rom_memory[38166] = 3'b110;
        rom_memory[38167] = 3'b110;
        rom_memory[38168] = 3'b110;
        rom_memory[38169] = 3'b111;
        rom_memory[38170] = 3'b111;
        rom_memory[38171] = 3'b111;
        rom_memory[38172] = 3'b111;
        rom_memory[38173] = 3'b111;
        rom_memory[38174] = 3'b111;
        rom_memory[38175] = 3'b111;
        rom_memory[38176] = 3'b111;
        rom_memory[38177] = 3'b111;
        rom_memory[38178] = 3'b111;
        rom_memory[38179] = 3'b111;
        rom_memory[38180] = 3'b111;
        rom_memory[38181] = 3'b111;
        rom_memory[38182] = 3'b111;
        rom_memory[38183] = 3'b111;
        rom_memory[38184] = 3'b111;
        rom_memory[38185] = 3'b110;
        rom_memory[38186] = 3'b110;
        rom_memory[38187] = 3'b110;
        rom_memory[38188] = 3'b110;
        rom_memory[38189] = 3'b110;
        rom_memory[38190] = 3'b110;
        rom_memory[38191] = 3'b110;
        rom_memory[38192] = 3'b110;
        rom_memory[38193] = 3'b110;
        rom_memory[38194] = 3'b110;
        rom_memory[38195] = 3'b110;
        rom_memory[38196] = 3'b110;
        rom_memory[38197] = 3'b110;
        rom_memory[38198] = 3'b110;
        rom_memory[38199] = 3'b110;
        rom_memory[38200] = 3'b110;
        rom_memory[38201] = 3'b110;
        rom_memory[38202] = 3'b110;
        rom_memory[38203] = 3'b111;
        rom_memory[38204] = 3'b111;
        rom_memory[38205] = 3'b111;
        rom_memory[38206] = 3'b111;
        rom_memory[38207] = 3'b111;
        rom_memory[38208] = 3'b111;
        rom_memory[38209] = 3'b111;
        rom_memory[38210] = 3'b111;
        rom_memory[38211] = 3'b111;
        rom_memory[38212] = 3'b111;
        rom_memory[38213] = 3'b111;
        rom_memory[38214] = 3'b111;
        rom_memory[38215] = 3'b111;
        rom_memory[38216] = 3'b111;
        rom_memory[38217] = 3'b110;
        rom_memory[38218] = 3'b111;
        rom_memory[38219] = 3'b111;
        rom_memory[38220] = 3'b111;
        rom_memory[38221] = 3'b110;
        rom_memory[38222] = 3'b111;
        rom_memory[38223] = 3'b111;
        rom_memory[38224] = 3'b110;
        rom_memory[38225] = 3'b110;
        rom_memory[38226] = 3'b111;
        rom_memory[38227] = 3'b000;
        rom_memory[38228] = 3'b000;
        rom_memory[38229] = 3'b000;
        rom_memory[38230] = 3'b110;
        rom_memory[38231] = 3'b110;
        rom_memory[38232] = 3'b110;
        rom_memory[38233] = 3'b110;
        rom_memory[38234] = 3'b110;
        rom_memory[38235] = 3'b110;
        rom_memory[38236] = 3'b110;
        rom_memory[38237] = 3'b110;
        rom_memory[38238] = 3'b110;
        rom_memory[38239] = 3'b111;
        rom_memory[38240] = 3'b111;
        rom_memory[38241] = 3'b000;
        rom_memory[38242] = 3'b000;
        rom_memory[38243] = 3'b111;
        rom_memory[38244] = 3'b111;
        rom_memory[38245] = 3'b100;
        rom_memory[38246] = 3'b000;
        rom_memory[38247] = 3'b000;
        rom_memory[38248] = 3'b110;
        rom_memory[38249] = 3'b111;
        rom_memory[38250] = 3'b111;
        rom_memory[38251] = 3'b111;
        rom_memory[38252] = 3'b111;
        rom_memory[38253] = 3'b111;
        rom_memory[38254] = 3'b111;
        rom_memory[38255] = 3'b011;
        rom_memory[38256] = 3'b011;
        rom_memory[38257] = 3'b111;
        rom_memory[38258] = 3'b111;
        rom_memory[38259] = 3'b111;
        rom_memory[38260] = 3'b111;
        rom_memory[38261] = 3'b110;
        rom_memory[38262] = 3'b110;
        rom_memory[38263] = 3'b110;
        rom_memory[38264] = 3'b110;
        rom_memory[38265] = 3'b110;
        rom_memory[38266] = 3'b110;
        rom_memory[38267] = 3'b110;
        rom_memory[38268] = 3'b110;
        rom_memory[38269] = 3'b110;
        rom_memory[38270] = 3'b110;
        rom_memory[38271] = 3'b110;
        rom_memory[38272] = 3'b110;
        rom_memory[38273] = 3'b110;
        rom_memory[38274] = 3'b110;
        rom_memory[38275] = 3'b110;
        rom_memory[38276] = 3'b110;
        rom_memory[38277] = 3'b110;
        rom_memory[38278] = 3'b110;
        rom_memory[38279] = 3'b110;
        rom_memory[38280] = 3'b110;
        rom_memory[38281] = 3'b110;
        rom_memory[38282] = 3'b110;
        rom_memory[38283] = 3'b110;
        rom_memory[38284] = 3'b110;
        rom_memory[38285] = 3'b110;
        rom_memory[38286] = 3'b110;
        rom_memory[38287] = 3'b110;
        rom_memory[38288] = 3'b110;
        rom_memory[38289] = 3'b110;
        rom_memory[38290] = 3'b110;
        rom_memory[38291] = 3'b110;
        rom_memory[38292] = 3'b110;
        rom_memory[38293] = 3'b110;
        rom_memory[38294] = 3'b110;
        rom_memory[38295] = 3'b110;
        rom_memory[38296] = 3'b110;
        rom_memory[38297] = 3'b110;
        rom_memory[38298] = 3'b110;
        rom_memory[38299] = 3'b110;
        rom_memory[38300] = 3'b110;
        rom_memory[38301] = 3'b110;
        rom_memory[38302] = 3'b110;
        rom_memory[38303] = 3'b110;
        rom_memory[38304] = 3'b110;
        rom_memory[38305] = 3'b110;
        rom_memory[38306] = 3'b110;
        rom_memory[38307] = 3'b110;
        rom_memory[38308] = 3'b110;
        rom_memory[38309] = 3'b110;
        rom_memory[38310] = 3'b110;
        rom_memory[38311] = 3'b110;
        rom_memory[38312] = 3'b110;
        rom_memory[38313] = 3'b110;
        rom_memory[38314] = 3'b110;
        rom_memory[38315] = 3'b110;
        rom_memory[38316] = 3'b110;
        rom_memory[38317] = 3'b110;
        rom_memory[38318] = 3'b111;
        rom_memory[38319] = 3'b110;
        rom_memory[38320] = 3'b000;
        rom_memory[38321] = 3'b000;
        rom_memory[38322] = 3'b000;
        rom_memory[38323] = 3'b000;
        rom_memory[38324] = 3'b000;
        rom_memory[38325] = 3'b110;
        rom_memory[38326] = 3'b000;
        rom_memory[38327] = 3'b000;
        rom_memory[38328] = 3'b000;
        rom_memory[38329] = 3'b000;
        rom_memory[38330] = 3'b000;
        rom_memory[38331] = 3'b000;
        rom_memory[38332] = 3'b000;
        rom_memory[38333] = 3'b000;
        rom_memory[38334] = 3'b100;
        rom_memory[38335] = 3'b111;
        rom_memory[38336] = 3'b111;
        rom_memory[38337] = 3'b110;
        rom_memory[38338] = 3'b110;
        rom_memory[38339] = 3'b110;
        rom_memory[38340] = 3'b110;
        rom_memory[38341] = 3'b110;
        rom_memory[38342] = 3'b110;
        rom_memory[38343] = 3'b110;
        rom_memory[38344] = 3'b110;
        rom_memory[38345] = 3'b110;
        rom_memory[38346] = 3'b110;
        rom_memory[38347] = 3'b110;
        rom_memory[38348] = 3'b110;
        rom_memory[38349] = 3'b110;
        rom_memory[38350] = 3'b110;
        rom_memory[38351] = 3'b110;
        rom_memory[38352] = 3'b110;
        rom_memory[38353] = 3'b110;
        rom_memory[38354] = 3'b110;
        rom_memory[38355] = 3'b110;
        rom_memory[38356] = 3'b110;
        rom_memory[38357] = 3'b110;
        rom_memory[38358] = 3'b110;
        rom_memory[38359] = 3'b110;
        rom_memory[38360] = 3'b110;
        rom_memory[38361] = 3'b110;
        rom_memory[38362] = 3'b110;
        rom_memory[38363] = 3'b110;
        rom_memory[38364] = 3'b110;
        rom_memory[38365] = 3'b111;
        rom_memory[38366] = 3'b111;
        rom_memory[38367] = 3'b111;
        rom_memory[38368] = 3'b111;
        rom_memory[38369] = 3'b111;
        rom_memory[38370] = 3'b111;
        rom_memory[38371] = 3'b111;
        rom_memory[38372] = 3'b111;
        rom_memory[38373] = 3'b111;
        rom_memory[38374] = 3'b111;
        rom_memory[38375] = 3'b111;
        rom_memory[38376] = 3'b111;
        rom_memory[38377] = 3'b111;
        rom_memory[38378] = 3'b111;
        rom_memory[38379] = 3'b111;
        rom_memory[38380] = 3'b111;
        rom_memory[38381] = 3'b111;
        rom_memory[38382] = 3'b111;
        rom_memory[38383] = 3'b111;
        rom_memory[38384] = 3'b111;
        rom_memory[38385] = 3'b111;
        rom_memory[38386] = 3'b111;
        rom_memory[38387] = 3'b111;
        rom_memory[38388] = 3'b111;
        rom_memory[38389] = 3'b111;
        rom_memory[38390] = 3'b111;
        rom_memory[38391] = 3'b111;
        rom_memory[38392] = 3'b111;
        rom_memory[38393] = 3'b111;
        rom_memory[38394] = 3'b111;
        rom_memory[38395] = 3'b111;
        rom_memory[38396] = 3'b111;
        rom_memory[38397] = 3'b111;
        rom_memory[38398] = 3'b111;
        rom_memory[38399] = 3'b111;
        rom_memory[38400] = 3'b110;
        rom_memory[38401] = 3'b110;
        rom_memory[38402] = 3'b110;
        rom_memory[38403] = 3'b110;
        rom_memory[38404] = 3'b110;
        rom_memory[38405] = 3'b110;
        rom_memory[38406] = 3'b110;
        rom_memory[38407] = 3'b110;
        rom_memory[38408] = 3'b110;
        rom_memory[38409] = 3'b111;
        rom_memory[38410] = 3'b111;
        rom_memory[38411] = 3'b111;
        rom_memory[38412] = 3'b111;
        rom_memory[38413] = 3'b111;
        rom_memory[38414] = 3'b111;
        rom_memory[38415] = 3'b111;
        rom_memory[38416] = 3'b111;
        rom_memory[38417] = 3'b111;
        rom_memory[38418] = 3'b111;
        rom_memory[38419] = 3'b111;
        rom_memory[38420] = 3'b111;
        rom_memory[38421] = 3'b111;
        rom_memory[38422] = 3'b111;
        rom_memory[38423] = 3'b111;
        rom_memory[38424] = 3'b110;
        rom_memory[38425] = 3'b110;
        rom_memory[38426] = 3'b110;
        rom_memory[38427] = 3'b110;
        rom_memory[38428] = 3'b110;
        rom_memory[38429] = 3'b110;
        rom_memory[38430] = 3'b110;
        rom_memory[38431] = 3'b110;
        rom_memory[38432] = 3'b110;
        rom_memory[38433] = 3'b110;
        rom_memory[38434] = 3'b110;
        rom_memory[38435] = 3'b110;
        rom_memory[38436] = 3'b110;
        rom_memory[38437] = 3'b110;
        rom_memory[38438] = 3'b110;
        rom_memory[38439] = 3'b110;
        rom_memory[38440] = 3'b110;
        rom_memory[38441] = 3'b110;
        rom_memory[38442] = 3'b110;
        rom_memory[38443] = 3'b111;
        rom_memory[38444] = 3'b111;
        rom_memory[38445] = 3'b111;
        rom_memory[38446] = 3'b111;
        rom_memory[38447] = 3'b111;
        rom_memory[38448] = 3'b111;
        rom_memory[38449] = 3'b111;
        rom_memory[38450] = 3'b111;
        rom_memory[38451] = 3'b111;
        rom_memory[38452] = 3'b110;
        rom_memory[38453] = 3'b110;
        rom_memory[38454] = 3'b110;
        rom_memory[38455] = 3'b110;
        rom_memory[38456] = 3'b110;
        rom_memory[38457] = 3'b100;
        rom_memory[38458] = 3'b100;
        rom_memory[38459] = 3'b110;
        rom_memory[38460] = 3'b100;
        rom_memory[38461] = 3'b110;
        rom_memory[38462] = 3'b111;
        rom_memory[38463] = 3'b110;
        rom_memory[38464] = 3'b110;
        rom_memory[38465] = 3'b110;
        rom_memory[38466] = 3'b110;
        rom_memory[38467] = 3'b000;
        rom_memory[38468] = 3'b000;
        rom_memory[38469] = 3'b000;
        rom_memory[38470] = 3'b110;
        rom_memory[38471] = 3'b110;
        rom_memory[38472] = 3'b110;
        rom_memory[38473] = 3'b110;
        rom_memory[38474] = 3'b110;
        rom_memory[38475] = 3'b110;
        rom_memory[38476] = 3'b111;
        rom_memory[38477] = 3'b110;
        rom_memory[38478] = 3'b000;
        rom_memory[38479] = 3'b111;
        rom_memory[38480] = 3'b100;
        rom_memory[38481] = 3'b000;
        rom_memory[38482] = 3'b000;
        rom_memory[38483] = 3'b000;
        rom_memory[38484] = 3'b110;
        rom_memory[38485] = 3'b000;
        rom_memory[38486] = 3'b000;
        rom_memory[38487] = 3'b000;
        rom_memory[38488] = 3'b111;
        rom_memory[38489] = 3'b111;
        rom_memory[38490] = 3'b111;
        rom_memory[38491] = 3'b111;
        rom_memory[38492] = 3'b111;
        rom_memory[38493] = 3'b111;
        rom_memory[38494] = 3'b111;
        rom_memory[38495] = 3'b111;
        rom_memory[38496] = 3'b011;
        rom_memory[38497] = 3'b111;
        rom_memory[38498] = 3'b111;
        rom_memory[38499] = 3'b111;
        rom_memory[38500] = 3'b111;
        rom_memory[38501] = 3'b111;
        rom_memory[38502] = 3'b110;
        rom_memory[38503] = 3'b110;
        rom_memory[38504] = 3'b110;
        rom_memory[38505] = 3'b110;
        rom_memory[38506] = 3'b110;
        rom_memory[38507] = 3'b110;
        rom_memory[38508] = 3'b110;
        rom_memory[38509] = 3'b110;
        rom_memory[38510] = 3'b110;
        rom_memory[38511] = 3'b110;
        rom_memory[38512] = 3'b110;
        rom_memory[38513] = 3'b110;
        rom_memory[38514] = 3'b110;
        rom_memory[38515] = 3'b110;
        rom_memory[38516] = 3'b110;
        rom_memory[38517] = 3'b110;
        rom_memory[38518] = 3'b110;
        rom_memory[38519] = 3'b110;
        rom_memory[38520] = 3'b110;
        rom_memory[38521] = 3'b110;
        rom_memory[38522] = 3'b110;
        rom_memory[38523] = 3'b110;
        rom_memory[38524] = 3'b110;
        rom_memory[38525] = 3'b110;
        rom_memory[38526] = 3'b110;
        rom_memory[38527] = 3'b110;
        rom_memory[38528] = 3'b110;
        rom_memory[38529] = 3'b110;
        rom_memory[38530] = 3'b110;
        rom_memory[38531] = 3'b110;
        rom_memory[38532] = 3'b110;
        rom_memory[38533] = 3'b110;
        rom_memory[38534] = 3'b110;
        rom_memory[38535] = 3'b110;
        rom_memory[38536] = 3'b110;
        rom_memory[38537] = 3'b110;
        rom_memory[38538] = 3'b110;
        rom_memory[38539] = 3'b110;
        rom_memory[38540] = 3'b110;
        rom_memory[38541] = 3'b110;
        rom_memory[38542] = 3'b110;
        rom_memory[38543] = 3'b110;
        rom_memory[38544] = 3'b110;
        rom_memory[38545] = 3'b110;
        rom_memory[38546] = 3'b110;
        rom_memory[38547] = 3'b110;
        rom_memory[38548] = 3'b110;
        rom_memory[38549] = 3'b110;
        rom_memory[38550] = 3'b110;
        rom_memory[38551] = 3'b110;
        rom_memory[38552] = 3'b110;
        rom_memory[38553] = 3'b110;
        rom_memory[38554] = 3'b110;
        rom_memory[38555] = 3'b110;
        rom_memory[38556] = 3'b110;
        rom_memory[38557] = 3'b110;
        rom_memory[38558] = 3'b110;
        rom_memory[38559] = 3'b111;
        rom_memory[38560] = 3'b110;
        rom_memory[38561] = 3'b000;
        rom_memory[38562] = 3'b000;
        rom_memory[38563] = 3'b000;
        rom_memory[38564] = 3'b000;
        rom_memory[38565] = 3'b000;
        rom_memory[38566] = 3'b110;
        rom_memory[38567] = 3'b000;
        rom_memory[38568] = 3'b000;
        rom_memory[38569] = 3'b000;
        rom_memory[38570] = 3'b000;
        rom_memory[38571] = 3'b000;
        rom_memory[38572] = 3'b000;
        rom_memory[38573] = 3'b000;
        rom_memory[38574] = 3'b000;
        rom_memory[38575] = 3'b000;
        rom_memory[38576] = 3'b111;
        rom_memory[38577] = 3'b111;
        rom_memory[38578] = 3'b110;
        rom_memory[38579] = 3'b110;
        rom_memory[38580] = 3'b110;
        rom_memory[38581] = 3'b110;
        rom_memory[38582] = 3'b110;
        rom_memory[38583] = 3'b110;
        rom_memory[38584] = 3'b110;
        rom_memory[38585] = 3'b110;
        rom_memory[38586] = 3'b110;
        rom_memory[38587] = 3'b110;
        rom_memory[38588] = 3'b110;
        rom_memory[38589] = 3'b110;
        rom_memory[38590] = 3'b110;
        rom_memory[38591] = 3'b110;
        rom_memory[38592] = 3'b110;
        rom_memory[38593] = 3'b110;
        rom_memory[38594] = 3'b110;
        rom_memory[38595] = 3'b110;
        rom_memory[38596] = 3'b110;
        rom_memory[38597] = 3'b110;
        rom_memory[38598] = 3'b110;
        rom_memory[38599] = 3'b110;
        rom_memory[38600] = 3'b110;
        rom_memory[38601] = 3'b110;
        rom_memory[38602] = 3'b110;
        rom_memory[38603] = 3'b110;
        rom_memory[38604] = 3'b110;
        rom_memory[38605] = 3'b110;
        rom_memory[38606] = 3'b111;
        rom_memory[38607] = 3'b111;
        rom_memory[38608] = 3'b111;
        rom_memory[38609] = 3'b111;
        rom_memory[38610] = 3'b111;
        rom_memory[38611] = 3'b111;
        rom_memory[38612] = 3'b111;
        rom_memory[38613] = 3'b111;
        rom_memory[38614] = 3'b111;
        rom_memory[38615] = 3'b111;
        rom_memory[38616] = 3'b111;
        rom_memory[38617] = 3'b111;
        rom_memory[38618] = 3'b111;
        rom_memory[38619] = 3'b111;
        rom_memory[38620] = 3'b111;
        rom_memory[38621] = 3'b111;
        rom_memory[38622] = 3'b111;
        rom_memory[38623] = 3'b111;
        rom_memory[38624] = 3'b111;
        rom_memory[38625] = 3'b111;
        rom_memory[38626] = 3'b111;
        rom_memory[38627] = 3'b111;
        rom_memory[38628] = 3'b111;
        rom_memory[38629] = 3'b111;
        rom_memory[38630] = 3'b111;
        rom_memory[38631] = 3'b111;
        rom_memory[38632] = 3'b111;
        rom_memory[38633] = 3'b111;
        rom_memory[38634] = 3'b111;
        rom_memory[38635] = 3'b111;
        rom_memory[38636] = 3'b111;
        rom_memory[38637] = 3'b111;
        rom_memory[38638] = 3'b111;
        rom_memory[38639] = 3'b111;
        rom_memory[38640] = 3'b110;
        rom_memory[38641] = 3'b110;
        rom_memory[38642] = 3'b110;
        rom_memory[38643] = 3'b110;
        rom_memory[38644] = 3'b110;
        rom_memory[38645] = 3'b110;
        rom_memory[38646] = 3'b110;
        rom_memory[38647] = 3'b110;
        rom_memory[38648] = 3'b110;
        rom_memory[38649] = 3'b111;
        rom_memory[38650] = 3'b111;
        rom_memory[38651] = 3'b111;
        rom_memory[38652] = 3'b111;
        rom_memory[38653] = 3'b111;
        rom_memory[38654] = 3'b111;
        rom_memory[38655] = 3'b111;
        rom_memory[38656] = 3'b111;
        rom_memory[38657] = 3'b111;
        rom_memory[38658] = 3'b111;
        rom_memory[38659] = 3'b111;
        rom_memory[38660] = 3'b111;
        rom_memory[38661] = 3'b111;
        rom_memory[38662] = 3'b111;
        rom_memory[38663] = 3'b111;
        rom_memory[38664] = 3'b110;
        rom_memory[38665] = 3'b110;
        rom_memory[38666] = 3'b110;
        rom_memory[38667] = 3'b110;
        rom_memory[38668] = 3'b110;
        rom_memory[38669] = 3'b110;
        rom_memory[38670] = 3'b110;
        rom_memory[38671] = 3'b110;
        rom_memory[38672] = 3'b110;
        rom_memory[38673] = 3'b110;
        rom_memory[38674] = 3'b110;
        rom_memory[38675] = 3'b110;
        rom_memory[38676] = 3'b110;
        rom_memory[38677] = 3'b110;
        rom_memory[38678] = 3'b110;
        rom_memory[38679] = 3'b110;
        rom_memory[38680] = 3'b110;
        rom_memory[38681] = 3'b110;
        rom_memory[38682] = 3'b110;
        rom_memory[38683] = 3'b111;
        rom_memory[38684] = 3'b111;
        rom_memory[38685] = 3'b111;
        rom_memory[38686] = 3'b111;
        rom_memory[38687] = 3'b111;
        rom_memory[38688] = 3'b111;
        rom_memory[38689] = 3'b111;
        rom_memory[38690] = 3'b111;
        rom_memory[38691] = 3'b111;
        rom_memory[38692] = 3'b110;
        rom_memory[38693] = 3'b110;
        rom_memory[38694] = 3'b111;
        rom_memory[38695] = 3'b110;
        rom_memory[38696] = 3'b110;
        rom_memory[38697] = 3'b000;
        rom_memory[38698] = 3'b000;
        rom_memory[38699] = 3'b100;
        rom_memory[38700] = 3'b100;
        rom_memory[38701] = 3'b110;
        rom_memory[38702] = 3'b111;
        rom_memory[38703] = 3'b110;
        rom_memory[38704] = 3'b110;
        rom_memory[38705] = 3'b110;
        rom_memory[38706] = 3'b110;
        rom_memory[38707] = 3'b100;
        rom_memory[38708] = 3'b110;
        rom_memory[38709] = 3'b110;
        rom_memory[38710] = 3'b110;
        rom_memory[38711] = 3'b110;
        rom_memory[38712] = 3'b110;
        rom_memory[38713] = 3'b110;
        rom_memory[38714] = 3'b110;
        rom_memory[38715] = 3'b110;
        rom_memory[38716] = 3'b111;
        rom_memory[38717] = 3'b100;
        rom_memory[38718] = 3'b000;
        rom_memory[38719] = 3'b110;
        rom_memory[38720] = 3'b100;
        rom_memory[38721] = 3'b000;
        rom_memory[38722] = 3'b000;
        rom_memory[38723] = 3'b110;
        rom_memory[38724] = 3'b100;
        rom_memory[38725] = 3'b110;
        rom_memory[38726] = 3'b110;
        rom_memory[38727] = 3'b110;
        rom_memory[38728] = 3'b111;
        rom_memory[38729] = 3'b110;
        rom_memory[38730] = 3'b110;
        rom_memory[38731] = 3'b110;
        rom_memory[38732] = 3'b111;
        rom_memory[38733] = 3'b111;
        rom_memory[38734] = 3'b111;
        rom_memory[38735] = 3'b111;
        rom_memory[38736] = 3'b111;
        rom_memory[38737] = 3'b111;
        rom_memory[38738] = 3'b111;
        rom_memory[38739] = 3'b111;
        rom_memory[38740] = 3'b111;
        rom_memory[38741] = 3'b111;
        rom_memory[38742] = 3'b110;
        rom_memory[38743] = 3'b110;
        rom_memory[38744] = 3'b110;
        rom_memory[38745] = 3'b110;
        rom_memory[38746] = 3'b110;
        rom_memory[38747] = 3'b110;
        rom_memory[38748] = 3'b110;
        rom_memory[38749] = 3'b110;
        rom_memory[38750] = 3'b110;
        rom_memory[38751] = 3'b110;
        rom_memory[38752] = 3'b110;
        rom_memory[38753] = 3'b110;
        rom_memory[38754] = 3'b110;
        rom_memory[38755] = 3'b110;
        rom_memory[38756] = 3'b110;
        rom_memory[38757] = 3'b110;
        rom_memory[38758] = 3'b110;
        rom_memory[38759] = 3'b110;
        rom_memory[38760] = 3'b110;
        rom_memory[38761] = 3'b110;
        rom_memory[38762] = 3'b110;
        rom_memory[38763] = 3'b110;
        rom_memory[38764] = 3'b110;
        rom_memory[38765] = 3'b110;
        rom_memory[38766] = 3'b110;
        rom_memory[38767] = 3'b110;
        rom_memory[38768] = 3'b110;
        rom_memory[38769] = 3'b110;
        rom_memory[38770] = 3'b110;
        rom_memory[38771] = 3'b110;
        rom_memory[38772] = 3'b110;
        rom_memory[38773] = 3'b110;
        rom_memory[38774] = 3'b110;
        rom_memory[38775] = 3'b110;
        rom_memory[38776] = 3'b110;
        rom_memory[38777] = 3'b110;
        rom_memory[38778] = 3'b110;
        rom_memory[38779] = 3'b110;
        rom_memory[38780] = 3'b110;
        rom_memory[38781] = 3'b110;
        rom_memory[38782] = 3'b110;
        rom_memory[38783] = 3'b110;
        rom_memory[38784] = 3'b110;
        rom_memory[38785] = 3'b110;
        rom_memory[38786] = 3'b110;
        rom_memory[38787] = 3'b110;
        rom_memory[38788] = 3'b110;
        rom_memory[38789] = 3'b110;
        rom_memory[38790] = 3'b110;
        rom_memory[38791] = 3'b110;
        rom_memory[38792] = 3'b110;
        rom_memory[38793] = 3'b110;
        rom_memory[38794] = 3'b110;
        rom_memory[38795] = 3'b110;
        rom_memory[38796] = 3'b110;
        rom_memory[38797] = 3'b110;
        rom_memory[38798] = 3'b110;
        rom_memory[38799] = 3'b110;
        rom_memory[38800] = 3'b111;
        rom_memory[38801] = 3'b110;
        rom_memory[38802] = 3'b000;
        rom_memory[38803] = 3'b000;
        rom_memory[38804] = 3'b000;
        rom_memory[38805] = 3'b000;
        rom_memory[38806] = 3'b000;
        rom_memory[38807] = 3'b110;
        rom_memory[38808] = 3'b000;
        rom_memory[38809] = 3'b000;
        rom_memory[38810] = 3'b000;
        rom_memory[38811] = 3'b000;
        rom_memory[38812] = 3'b000;
        rom_memory[38813] = 3'b000;
        rom_memory[38814] = 3'b000;
        rom_memory[38815] = 3'b000;
        rom_memory[38816] = 3'b000;
        rom_memory[38817] = 3'b110;
        rom_memory[38818] = 3'b111;
        rom_memory[38819] = 3'b110;
        rom_memory[38820] = 3'b110;
        rom_memory[38821] = 3'b110;
        rom_memory[38822] = 3'b110;
        rom_memory[38823] = 3'b110;
        rom_memory[38824] = 3'b110;
        rom_memory[38825] = 3'b110;
        rom_memory[38826] = 3'b110;
        rom_memory[38827] = 3'b110;
        rom_memory[38828] = 3'b110;
        rom_memory[38829] = 3'b110;
        rom_memory[38830] = 3'b110;
        rom_memory[38831] = 3'b110;
        rom_memory[38832] = 3'b110;
        rom_memory[38833] = 3'b110;
        rom_memory[38834] = 3'b110;
        rom_memory[38835] = 3'b110;
        rom_memory[38836] = 3'b110;
        rom_memory[38837] = 3'b110;
        rom_memory[38838] = 3'b110;
        rom_memory[38839] = 3'b110;
        rom_memory[38840] = 3'b110;
        rom_memory[38841] = 3'b110;
        rom_memory[38842] = 3'b110;
        rom_memory[38843] = 3'b110;
        rom_memory[38844] = 3'b110;
        rom_memory[38845] = 3'b110;
        rom_memory[38846] = 3'b111;
        rom_memory[38847] = 3'b111;
        rom_memory[38848] = 3'b111;
        rom_memory[38849] = 3'b111;
        rom_memory[38850] = 3'b111;
        rom_memory[38851] = 3'b111;
        rom_memory[38852] = 3'b111;
        rom_memory[38853] = 3'b111;
        rom_memory[38854] = 3'b111;
        rom_memory[38855] = 3'b111;
        rom_memory[38856] = 3'b111;
        rom_memory[38857] = 3'b111;
        rom_memory[38858] = 3'b111;
        rom_memory[38859] = 3'b111;
        rom_memory[38860] = 3'b111;
        rom_memory[38861] = 3'b111;
        rom_memory[38862] = 3'b111;
        rom_memory[38863] = 3'b111;
        rom_memory[38864] = 3'b111;
        rom_memory[38865] = 3'b111;
        rom_memory[38866] = 3'b111;
        rom_memory[38867] = 3'b111;
        rom_memory[38868] = 3'b111;
        rom_memory[38869] = 3'b111;
        rom_memory[38870] = 3'b111;
        rom_memory[38871] = 3'b111;
        rom_memory[38872] = 3'b111;
        rom_memory[38873] = 3'b111;
        rom_memory[38874] = 3'b111;
        rom_memory[38875] = 3'b111;
        rom_memory[38876] = 3'b111;
        rom_memory[38877] = 3'b111;
        rom_memory[38878] = 3'b111;
        rom_memory[38879] = 3'b111;
        rom_memory[38880] = 3'b110;
        rom_memory[38881] = 3'b110;
        rom_memory[38882] = 3'b110;
        rom_memory[38883] = 3'b110;
        rom_memory[38884] = 3'b110;
        rom_memory[38885] = 3'b110;
        rom_memory[38886] = 3'b110;
        rom_memory[38887] = 3'b110;
        rom_memory[38888] = 3'b110;
        rom_memory[38889] = 3'b110;
        rom_memory[38890] = 3'b111;
        rom_memory[38891] = 3'b111;
        rom_memory[38892] = 3'b111;
        rom_memory[38893] = 3'b111;
        rom_memory[38894] = 3'b111;
        rom_memory[38895] = 3'b111;
        rom_memory[38896] = 3'b111;
        rom_memory[38897] = 3'b111;
        rom_memory[38898] = 3'b111;
        rom_memory[38899] = 3'b111;
        rom_memory[38900] = 3'b111;
        rom_memory[38901] = 3'b111;
        rom_memory[38902] = 3'b111;
        rom_memory[38903] = 3'b110;
        rom_memory[38904] = 3'b110;
        rom_memory[38905] = 3'b110;
        rom_memory[38906] = 3'b110;
        rom_memory[38907] = 3'b110;
        rom_memory[38908] = 3'b110;
        rom_memory[38909] = 3'b110;
        rom_memory[38910] = 3'b110;
        rom_memory[38911] = 3'b110;
        rom_memory[38912] = 3'b110;
        rom_memory[38913] = 3'b110;
        rom_memory[38914] = 3'b110;
        rom_memory[38915] = 3'b110;
        rom_memory[38916] = 3'b110;
        rom_memory[38917] = 3'b110;
        rom_memory[38918] = 3'b110;
        rom_memory[38919] = 3'b110;
        rom_memory[38920] = 3'b110;
        rom_memory[38921] = 3'b110;
        rom_memory[38922] = 3'b110;
        rom_memory[38923] = 3'b111;
        rom_memory[38924] = 3'b111;
        rom_memory[38925] = 3'b111;
        rom_memory[38926] = 3'b111;
        rom_memory[38927] = 3'b111;
        rom_memory[38928] = 3'b111;
        rom_memory[38929] = 3'b111;
        rom_memory[38930] = 3'b111;
        rom_memory[38931] = 3'b111;
        rom_memory[38932] = 3'b111;
        rom_memory[38933] = 3'b111;
        rom_memory[38934] = 3'b111;
        rom_memory[38935] = 3'b111;
        rom_memory[38936] = 3'b111;
        rom_memory[38937] = 3'b111;
        rom_memory[38938] = 3'b000;
        rom_memory[38939] = 3'b110;
        rom_memory[38940] = 3'b110;
        rom_memory[38941] = 3'b110;
        rom_memory[38942] = 3'b110;
        rom_memory[38943] = 3'b110;
        rom_memory[38944] = 3'b110;
        rom_memory[38945] = 3'b100;
        rom_memory[38946] = 3'b110;
        rom_memory[38947] = 3'b110;
        rom_memory[38948] = 3'b110;
        rom_memory[38949] = 3'b111;
        rom_memory[38950] = 3'b110;
        rom_memory[38951] = 3'b110;
        rom_memory[38952] = 3'b110;
        rom_memory[38953] = 3'b110;
        rom_memory[38954] = 3'b110;
        rom_memory[38955] = 3'b110;
        rom_memory[38956] = 3'b111;
        rom_memory[38957] = 3'b000;
        rom_memory[38958] = 3'b000;
        rom_memory[38959] = 3'b000;
        rom_memory[38960] = 3'b000;
        rom_memory[38961] = 3'b000;
        rom_memory[38962] = 3'b111;
        rom_memory[38963] = 3'b111;
        rom_memory[38964] = 3'b110;
        rom_memory[38965] = 3'b110;
        rom_memory[38966] = 3'b111;
        rom_memory[38967] = 3'b110;
        rom_memory[38968] = 3'b110;
        rom_memory[38969] = 3'b110;
        rom_memory[38970] = 3'b110;
        rom_memory[38971] = 3'b110;
        rom_memory[38972] = 3'b110;
        rom_memory[38973] = 3'b110;
        rom_memory[38974] = 3'b111;
        rom_memory[38975] = 3'b111;
        rom_memory[38976] = 3'b111;
        rom_memory[38977] = 3'b111;
        rom_memory[38978] = 3'b111;
        rom_memory[38979] = 3'b111;
        rom_memory[38980] = 3'b111;
        rom_memory[38981] = 3'b111;
        rom_memory[38982] = 3'b110;
        rom_memory[38983] = 3'b110;
        rom_memory[38984] = 3'b110;
        rom_memory[38985] = 3'b110;
        rom_memory[38986] = 3'b110;
        rom_memory[38987] = 3'b110;
        rom_memory[38988] = 3'b110;
        rom_memory[38989] = 3'b110;
        rom_memory[38990] = 3'b110;
        rom_memory[38991] = 3'b110;
        rom_memory[38992] = 3'b110;
        rom_memory[38993] = 3'b110;
        rom_memory[38994] = 3'b110;
        rom_memory[38995] = 3'b110;
        rom_memory[38996] = 3'b110;
        rom_memory[38997] = 3'b110;
        rom_memory[38998] = 3'b110;
        rom_memory[38999] = 3'b110;
        rom_memory[39000] = 3'b110;
        rom_memory[39001] = 3'b110;
        rom_memory[39002] = 3'b110;
        rom_memory[39003] = 3'b110;
        rom_memory[39004] = 3'b110;
        rom_memory[39005] = 3'b110;
        rom_memory[39006] = 3'b110;
        rom_memory[39007] = 3'b110;
        rom_memory[39008] = 3'b110;
        rom_memory[39009] = 3'b110;
        rom_memory[39010] = 3'b110;
        rom_memory[39011] = 3'b110;
        rom_memory[39012] = 3'b110;
        rom_memory[39013] = 3'b110;
        rom_memory[39014] = 3'b110;
        rom_memory[39015] = 3'b110;
        rom_memory[39016] = 3'b110;
        rom_memory[39017] = 3'b110;
        rom_memory[39018] = 3'b110;
        rom_memory[39019] = 3'b110;
        rom_memory[39020] = 3'b110;
        rom_memory[39021] = 3'b110;
        rom_memory[39022] = 3'b110;
        rom_memory[39023] = 3'b110;
        rom_memory[39024] = 3'b110;
        rom_memory[39025] = 3'b110;
        rom_memory[39026] = 3'b110;
        rom_memory[39027] = 3'b110;
        rom_memory[39028] = 3'b110;
        rom_memory[39029] = 3'b110;
        rom_memory[39030] = 3'b110;
        rom_memory[39031] = 3'b110;
        rom_memory[39032] = 3'b110;
        rom_memory[39033] = 3'b110;
        rom_memory[39034] = 3'b110;
        rom_memory[39035] = 3'b110;
        rom_memory[39036] = 3'b110;
        rom_memory[39037] = 3'b110;
        rom_memory[39038] = 3'b110;
        rom_memory[39039] = 3'b110;
        rom_memory[39040] = 3'b110;
        rom_memory[39041] = 3'b111;
        rom_memory[39042] = 3'b110;
        rom_memory[39043] = 3'b000;
        rom_memory[39044] = 3'b000;
        rom_memory[39045] = 3'b000;
        rom_memory[39046] = 3'b000;
        rom_memory[39047] = 3'b000;
        rom_memory[39048] = 3'b110;
        rom_memory[39049] = 3'b000;
        rom_memory[39050] = 3'b000;
        rom_memory[39051] = 3'b000;
        rom_memory[39052] = 3'b000;
        rom_memory[39053] = 3'b000;
        rom_memory[39054] = 3'b000;
        rom_memory[39055] = 3'b000;
        rom_memory[39056] = 3'b000;
        rom_memory[39057] = 3'b000;
        rom_memory[39058] = 3'b110;
        rom_memory[39059] = 3'b111;
        rom_memory[39060] = 3'b110;
        rom_memory[39061] = 3'b110;
        rom_memory[39062] = 3'b110;
        rom_memory[39063] = 3'b110;
        rom_memory[39064] = 3'b110;
        rom_memory[39065] = 3'b110;
        rom_memory[39066] = 3'b110;
        rom_memory[39067] = 3'b110;
        rom_memory[39068] = 3'b110;
        rom_memory[39069] = 3'b110;
        rom_memory[39070] = 3'b110;
        rom_memory[39071] = 3'b110;
        rom_memory[39072] = 3'b110;
        rom_memory[39073] = 3'b110;
        rom_memory[39074] = 3'b110;
        rom_memory[39075] = 3'b110;
        rom_memory[39076] = 3'b110;
        rom_memory[39077] = 3'b110;
        rom_memory[39078] = 3'b110;
        rom_memory[39079] = 3'b110;
        rom_memory[39080] = 3'b110;
        rom_memory[39081] = 3'b110;
        rom_memory[39082] = 3'b110;
        rom_memory[39083] = 3'b110;
        rom_memory[39084] = 3'b110;
        rom_memory[39085] = 3'b110;
        rom_memory[39086] = 3'b110;
        rom_memory[39087] = 3'b110;
        rom_memory[39088] = 3'b110;
        rom_memory[39089] = 3'b111;
        rom_memory[39090] = 3'b111;
        rom_memory[39091] = 3'b111;
        rom_memory[39092] = 3'b111;
        rom_memory[39093] = 3'b111;
        rom_memory[39094] = 3'b111;
        rom_memory[39095] = 3'b111;
        rom_memory[39096] = 3'b111;
        rom_memory[39097] = 3'b111;
        rom_memory[39098] = 3'b111;
        rom_memory[39099] = 3'b111;
        rom_memory[39100] = 3'b111;
        rom_memory[39101] = 3'b111;
        rom_memory[39102] = 3'b111;
        rom_memory[39103] = 3'b111;
        rom_memory[39104] = 3'b111;
        rom_memory[39105] = 3'b111;
        rom_memory[39106] = 3'b111;
        rom_memory[39107] = 3'b111;
        rom_memory[39108] = 3'b111;
        rom_memory[39109] = 3'b111;
        rom_memory[39110] = 3'b111;
        rom_memory[39111] = 3'b111;
        rom_memory[39112] = 3'b111;
        rom_memory[39113] = 3'b111;
        rom_memory[39114] = 3'b111;
        rom_memory[39115] = 3'b111;
        rom_memory[39116] = 3'b111;
        rom_memory[39117] = 3'b111;
        rom_memory[39118] = 3'b111;
        rom_memory[39119] = 3'b111;
        rom_memory[39120] = 3'b110;
        rom_memory[39121] = 3'b110;
        rom_memory[39122] = 3'b110;
        rom_memory[39123] = 3'b110;
        rom_memory[39124] = 3'b110;
        rom_memory[39125] = 3'b110;
        rom_memory[39126] = 3'b110;
        rom_memory[39127] = 3'b110;
        rom_memory[39128] = 3'b110;
        rom_memory[39129] = 3'b110;
        rom_memory[39130] = 3'b111;
        rom_memory[39131] = 3'b111;
        rom_memory[39132] = 3'b111;
        rom_memory[39133] = 3'b111;
        rom_memory[39134] = 3'b111;
        rom_memory[39135] = 3'b111;
        rom_memory[39136] = 3'b111;
        rom_memory[39137] = 3'b111;
        rom_memory[39138] = 3'b111;
        rom_memory[39139] = 3'b111;
        rom_memory[39140] = 3'b111;
        rom_memory[39141] = 3'b111;
        rom_memory[39142] = 3'b111;
        rom_memory[39143] = 3'b110;
        rom_memory[39144] = 3'b110;
        rom_memory[39145] = 3'b110;
        rom_memory[39146] = 3'b110;
        rom_memory[39147] = 3'b110;
        rom_memory[39148] = 3'b110;
        rom_memory[39149] = 3'b110;
        rom_memory[39150] = 3'b110;
        rom_memory[39151] = 3'b110;
        rom_memory[39152] = 3'b110;
        rom_memory[39153] = 3'b110;
        rom_memory[39154] = 3'b110;
        rom_memory[39155] = 3'b110;
        rom_memory[39156] = 3'b110;
        rom_memory[39157] = 3'b110;
        rom_memory[39158] = 3'b110;
        rom_memory[39159] = 3'b110;
        rom_memory[39160] = 3'b110;
        rom_memory[39161] = 3'b110;
        rom_memory[39162] = 3'b111;
        rom_memory[39163] = 3'b111;
        rom_memory[39164] = 3'b111;
        rom_memory[39165] = 3'b111;
        rom_memory[39166] = 3'b111;
        rom_memory[39167] = 3'b111;
        rom_memory[39168] = 3'b111;
        rom_memory[39169] = 3'b111;
        rom_memory[39170] = 3'b111;
        rom_memory[39171] = 3'b111;
        rom_memory[39172] = 3'b111;
        rom_memory[39173] = 3'b111;
        rom_memory[39174] = 3'b111;
        rom_memory[39175] = 3'b111;
        rom_memory[39176] = 3'b010;
        rom_memory[39177] = 3'b000;
        rom_memory[39178] = 3'b000;
        rom_memory[39179] = 3'b000;
        rom_memory[39180] = 3'b000;
        rom_memory[39181] = 3'b110;
        rom_memory[39182] = 3'b110;
        rom_memory[39183] = 3'b110;
        rom_memory[39184] = 3'b100;
        rom_memory[39185] = 3'b100;
        rom_memory[39186] = 3'b100;
        rom_memory[39187] = 3'b100;
        rom_memory[39188] = 3'b111;
        rom_memory[39189] = 3'b111;
        rom_memory[39190] = 3'b111;
        rom_memory[39191] = 3'b110;
        rom_memory[39192] = 3'b110;
        rom_memory[39193] = 3'b110;
        rom_memory[39194] = 3'b110;
        rom_memory[39195] = 3'b110;
        rom_memory[39196] = 3'b111;
        rom_memory[39197] = 3'b000;
        rom_memory[39198] = 3'b000;
        rom_memory[39199] = 3'b100;
        rom_memory[39200] = 3'b000;
        rom_memory[39201] = 3'b000;
        rom_memory[39202] = 3'b110;
        rom_memory[39203] = 3'b111;
        rom_memory[39204] = 3'b110;
        rom_memory[39205] = 3'b110;
        rom_memory[39206] = 3'b110;
        rom_memory[39207] = 3'b110;
        rom_memory[39208] = 3'b110;
        rom_memory[39209] = 3'b110;
        rom_memory[39210] = 3'b110;
        rom_memory[39211] = 3'b110;
        rom_memory[39212] = 3'b110;
        rom_memory[39213] = 3'b110;
        rom_memory[39214] = 3'b110;
        rom_memory[39215] = 3'b111;
        rom_memory[39216] = 3'b111;
        rom_memory[39217] = 3'b111;
        rom_memory[39218] = 3'b111;
        rom_memory[39219] = 3'b111;
        rom_memory[39220] = 3'b111;
        rom_memory[39221] = 3'b111;
        rom_memory[39222] = 3'b110;
        rom_memory[39223] = 3'b110;
        rom_memory[39224] = 3'b110;
        rom_memory[39225] = 3'b110;
        rom_memory[39226] = 3'b110;
        rom_memory[39227] = 3'b110;
        rom_memory[39228] = 3'b110;
        rom_memory[39229] = 3'b110;
        rom_memory[39230] = 3'b110;
        rom_memory[39231] = 3'b110;
        rom_memory[39232] = 3'b110;
        rom_memory[39233] = 3'b110;
        rom_memory[39234] = 3'b110;
        rom_memory[39235] = 3'b110;
        rom_memory[39236] = 3'b110;
        rom_memory[39237] = 3'b110;
        rom_memory[39238] = 3'b110;
        rom_memory[39239] = 3'b110;
        rom_memory[39240] = 3'b110;
        rom_memory[39241] = 3'b110;
        rom_memory[39242] = 3'b110;
        rom_memory[39243] = 3'b110;
        rom_memory[39244] = 3'b110;
        rom_memory[39245] = 3'b110;
        rom_memory[39246] = 3'b110;
        rom_memory[39247] = 3'b110;
        rom_memory[39248] = 3'b110;
        rom_memory[39249] = 3'b110;
        rom_memory[39250] = 3'b110;
        rom_memory[39251] = 3'b110;
        rom_memory[39252] = 3'b110;
        rom_memory[39253] = 3'b110;
        rom_memory[39254] = 3'b110;
        rom_memory[39255] = 3'b110;
        rom_memory[39256] = 3'b110;
        rom_memory[39257] = 3'b110;
        rom_memory[39258] = 3'b110;
        rom_memory[39259] = 3'b110;
        rom_memory[39260] = 3'b110;
        rom_memory[39261] = 3'b110;
        rom_memory[39262] = 3'b110;
        rom_memory[39263] = 3'b110;
        rom_memory[39264] = 3'b110;
        rom_memory[39265] = 3'b110;
        rom_memory[39266] = 3'b110;
        rom_memory[39267] = 3'b110;
        rom_memory[39268] = 3'b110;
        rom_memory[39269] = 3'b110;
        rom_memory[39270] = 3'b110;
        rom_memory[39271] = 3'b110;
        rom_memory[39272] = 3'b110;
        rom_memory[39273] = 3'b110;
        rom_memory[39274] = 3'b110;
        rom_memory[39275] = 3'b110;
        rom_memory[39276] = 3'b110;
        rom_memory[39277] = 3'b110;
        rom_memory[39278] = 3'b110;
        rom_memory[39279] = 3'b110;
        rom_memory[39280] = 3'b110;
        rom_memory[39281] = 3'b110;
        rom_memory[39282] = 3'b111;
        rom_memory[39283] = 3'b110;
        rom_memory[39284] = 3'b000;
        rom_memory[39285] = 3'b000;
        rom_memory[39286] = 3'b000;
        rom_memory[39287] = 3'b000;
        rom_memory[39288] = 3'b000;
        rom_memory[39289] = 3'b000;
        rom_memory[39290] = 3'b000;
        rom_memory[39291] = 3'b000;
        rom_memory[39292] = 3'b000;
        rom_memory[39293] = 3'b000;
        rom_memory[39294] = 3'b000;
        rom_memory[39295] = 3'b000;
        rom_memory[39296] = 3'b000;
        rom_memory[39297] = 3'b000;
        rom_memory[39298] = 3'b000;
        rom_memory[39299] = 3'b110;
        rom_memory[39300] = 3'b111;
        rom_memory[39301] = 3'b111;
        rom_memory[39302] = 3'b110;
        rom_memory[39303] = 3'b110;
        rom_memory[39304] = 3'b110;
        rom_memory[39305] = 3'b110;
        rom_memory[39306] = 3'b110;
        rom_memory[39307] = 3'b110;
        rom_memory[39308] = 3'b110;
        rom_memory[39309] = 3'b110;
        rom_memory[39310] = 3'b110;
        rom_memory[39311] = 3'b110;
        rom_memory[39312] = 3'b110;
        rom_memory[39313] = 3'b110;
        rom_memory[39314] = 3'b110;
        rom_memory[39315] = 3'b110;
        rom_memory[39316] = 3'b110;
        rom_memory[39317] = 3'b110;
        rom_memory[39318] = 3'b110;
        rom_memory[39319] = 3'b110;
        rom_memory[39320] = 3'b110;
        rom_memory[39321] = 3'b110;
        rom_memory[39322] = 3'b110;
        rom_memory[39323] = 3'b110;
        rom_memory[39324] = 3'b110;
        rom_memory[39325] = 3'b110;
        rom_memory[39326] = 3'b110;
        rom_memory[39327] = 3'b110;
        rom_memory[39328] = 3'b111;
        rom_memory[39329] = 3'b110;
        rom_memory[39330] = 3'b111;
        rom_memory[39331] = 3'b111;
        rom_memory[39332] = 3'b111;
        rom_memory[39333] = 3'b111;
        rom_memory[39334] = 3'b111;
        rom_memory[39335] = 3'b111;
        rom_memory[39336] = 3'b111;
        rom_memory[39337] = 3'b111;
        rom_memory[39338] = 3'b111;
        rom_memory[39339] = 3'b111;
        rom_memory[39340] = 3'b111;
        rom_memory[39341] = 3'b111;
        rom_memory[39342] = 3'b111;
        rom_memory[39343] = 3'b111;
        rom_memory[39344] = 3'b111;
        rom_memory[39345] = 3'b111;
        rom_memory[39346] = 3'b111;
        rom_memory[39347] = 3'b111;
        rom_memory[39348] = 3'b111;
        rom_memory[39349] = 3'b111;
        rom_memory[39350] = 3'b111;
        rom_memory[39351] = 3'b111;
        rom_memory[39352] = 3'b111;
        rom_memory[39353] = 3'b111;
        rom_memory[39354] = 3'b111;
        rom_memory[39355] = 3'b111;
        rom_memory[39356] = 3'b111;
        rom_memory[39357] = 3'b111;
        rom_memory[39358] = 3'b111;
        rom_memory[39359] = 3'b111;
        rom_memory[39360] = 3'b110;
        rom_memory[39361] = 3'b110;
        rom_memory[39362] = 3'b110;
        rom_memory[39363] = 3'b110;
        rom_memory[39364] = 3'b110;
        rom_memory[39365] = 3'b110;
        rom_memory[39366] = 3'b110;
        rom_memory[39367] = 3'b110;
        rom_memory[39368] = 3'b110;
        rom_memory[39369] = 3'b110;
        rom_memory[39370] = 3'b111;
        rom_memory[39371] = 3'b111;
        rom_memory[39372] = 3'b111;
        rom_memory[39373] = 3'b111;
        rom_memory[39374] = 3'b111;
        rom_memory[39375] = 3'b111;
        rom_memory[39376] = 3'b111;
        rom_memory[39377] = 3'b111;
        rom_memory[39378] = 3'b111;
        rom_memory[39379] = 3'b111;
        rom_memory[39380] = 3'b111;
        rom_memory[39381] = 3'b110;
        rom_memory[39382] = 3'b110;
        rom_memory[39383] = 3'b110;
        rom_memory[39384] = 3'b110;
        rom_memory[39385] = 3'b110;
        rom_memory[39386] = 3'b110;
        rom_memory[39387] = 3'b110;
        rom_memory[39388] = 3'b110;
        rom_memory[39389] = 3'b110;
        rom_memory[39390] = 3'b110;
        rom_memory[39391] = 3'b110;
        rom_memory[39392] = 3'b110;
        rom_memory[39393] = 3'b110;
        rom_memory[39394] = 3'b110;
        rom_memory[39395] = 3'b110;
        rom_memory[39396] = 3'b110;
        rom_memory[39397] = 3'b110;
        rom_memory[39398] = 3'b110;
        rom_memory[39399] = 3'b110;
        rom_memory[39400] = 3'b110;
        rom_memory[39401] = 3'b110;
        rom_memory[39402] = 3'b111;
        rom_memory[39403] = 3'b111;
        rom_memory[39404] = 3'b111;
        rom_memory[39405] = 3'b111;
        rom_memory[39406] = 3'b111;
        rom_memory[39407] = 3'b111;
        rom_memory[39408] = 3'b111;
        rom_memory[39409] = 3'b111;
        rom_memory[39410] = 3'b111;
        rom_memory[39411] = 3'b111;
        rom_memory[39412] = 3'b111;
        rom_memory[39413] = 3'b111;
        rom_memory[39414] = 3'b111;
        rom_memory[39415] = 3'b010;
        rom_memory[39416] = 3'b000;
        rom_memory[39417] = 3'b000;
        rom_memory[39418] = 3'b000;
        rom_memory[39419] = 3'b000;
        rom_memory[39420] = 3'b000;
        rom_memory[39421] = 3'b110;
        rom_memory[39422] = 3'b100;
        rom_memory[39423] = 3'b100;
        rom_memory[39424] = 3'b100;
        rom_memory[39425] = 3'b111;
        rom_memory[39426] = 3'b111;
        rom_memory[39427] = 3'b111;
        rom_memory[39428] = 3'b111;
        rom_memory[39429] = 3'b111;
        rom_memory[39430] = 3'b111;
        rom_memory[39431] = 3'b110;
        rom_memory[39432] = 3'b110;
        rom_memory[39433] = 3'b110;
        rom_memory[39434] = 3'b110;
        rom_memory[39435] = 3'b110;
        rom_memory[39436] = 3'b110;
        rom_memory[39437] = 3'b000;
        rom_memory[39438] = 3'b000;
        rom_memory[39439] = 3'b111;
        rom_memory[39440] = 3'b100;
        rom_memory[39441] = 3'b100;
        rom_memory[39442] = 3'b111;
        rom_memory[39443] = 3'b111;
        rom_memory[39444] = 3'b110;
        rom_memory[39445] = 3'b110;
        rom_memory[39446] = 3'b110;
        rom_memory[39447] = 3'b110;
        rom_memory[39448] = 3'b110;
        rom_memory[39449] = 3'b110;
        rom_memory[39450] = 3'b110;
        rom_memory[39451] = 3'b110;
        rom_memory[39452] = 3'b110;
        rom_memory[39453] = 3'b110;
        rom_memory[39454] = 3'b110;
        rom_memory[39455] = 3'b110;
        rom_memory[39456] = 3'b111;
        rom_memory[39457] = 3'b111;
        rom_memory[39458] = 3'b111;
        rom_memory[39459] = 3'b111;
        rom_memory[39460] = 3'b111;
        rom_memory[39461] = 3'b111;
        rom_memory[39462] = 3'b110;
        rom_memory[39463] = 3'b110;
        rom_memory[39464] = 3'b110;
        rom_memory[39465] = 3'b110;
        rom_memory[39466] = 3'b110;
        rom_memory[39467] = 3'b110;
        rom_memory[39468] = 3'b110;
        rom_memory[39469] = 3'b110;
        rom_memory[39470] = 3'b110;
        rom_memory[39471] = 3'b110;
        rom_memory[39472] = 3'b110;
        rom_memory[39473] = 3'b110;
        rom_memory[39474] = 3'b110;
        rom_memory[39475] = 3'b110;
        rom_memory[39476] = 3'b110;
        rom_memory[39477] = 3'b110;
        rom_memory[39478] = 3'b110;
        rom_memory[39479] = 3'b110;
        rom_memory[39480] = 3'b110;
        rom_memory[39481] = 3'b110;
        rom_memory[39482] = 3'b110;
        rom_memory[39483] = 3'b110;
        rom_memory[39484] = 3'b110;
        rom_memory[39485] = 3'b110;
        rom_memory[39486] = 3'b110;
        rom_memory[39487] = 3'b110;
        rom_memory[39488] = 3'b110;
        rom_memory[39489] = 3'b110;
        rom_memory[39490] = 3'b110;
        rom_memory[39491] = 3'b110;
        rom_memory[39492] = 3'b110;
        rom_memory[39493] = 3'b110;
        rom_memory[39494] = 3'b110;
        rom_memory[39495] = 3'b110;
        rom_memory[39496] = 3'b110;
        rom_memory[39497] = 3'b110;
        rom_memory[39498] = 3'b110;
        rom_memory[39499] = 3'b110;
        rom_memory[39500] = 3'b110;
        rom_memory[39501] = 3'b110;
        rom_memory[39502] = 3'b110;
        rom_memory[39503] = 3'b110;
        rom_memory[39504] = 3'b110;
        rom_memory[39505] = 3'b110;
        rom_memory[39506] = 3'b110;
        rom_memory[39507] = 3'b110;
        rom_memory[39508] = 3'b110;
        rom_memory[39509] = 3'b110;
        rom_memory[39510] = 3'b110;
        rom_memory[39511] = 3'b110;
        rom_memory[39512] = 3'b110;
        rom_memory[39513] = 3'b110;
        rom_memory[39514] = 3'b110;
        rom_memory[39515] = 3'b110;
        rom_memory[39516] = 3'b110;
        rom_memory[39517] = 3'b110;
        rom_memory[39518] = 3'b110;
        rom_memory[39519] = 3'b110;
        rom_memory[39520] = 3'b110;
        rom_memory[39521] = 3'b110;
        rom_memory[39522] = 3'b110;
        rom_memory[39523] = 3'b110;
        rom_memory[39524] = 3'b110;
        rom_memory[39525] = 3'b000;
        rom_memory[39526] = 3'b000;
        rom_memory[39527] = 3'b000;
        rom_memory[39528] = 3'b000;
        rom_memory[39529] = 3'b000;
        rom_memory[39530] = 3'b000;
        rom_memory[39531] = 3'b000;
        rom_memory[39532] = 3'b000;
        rom_memory[39533] = 3'b000;
        rom_memory[39534] = 3'b000;
        rom_memory[39535] = 3'b000;
        rom_memory[39536] = 3'b000;
        rom_memory[39537] = 3'b000;
        rom_memory[39538] = 3'b000;
        rom_memory[39539] = 3'b000;
        rom_memory[39540] = 3'b000;
        rom_memory[39541] = 3'b111;
        rom_memory[39542] = 3'b111;
        rom_memory[39543] = 3'b110;
        rom_memory[39544] = 3'b110;
        rom_memory[39545] = 3'b110;
        rom_memory[39546] = 3'b110;
        rom_memory[39547] = 3'b110;
        rom_memory[39548] = 3'b110;
        rom_memory[39549] = 3'b110;
        rom_memory[39550] = 3'b110;
        rom_memory[39551] = 3'b110;
        rom_memory[39552] = 3'b110;
        rom_memory[39553] = 3'b110;
        rom_memory[39554] = 3'b110;
        rom_memory[39555] = 3'b110;
        rom_memory[39556] = 3'b110;
        rom_memory[39557] = 3'b110;
        rom_memory[39558] = 3'b110;
        rom_memory[39559] = 3'b110;
        rom_memory[39560] = 3'b110;
        rom_memory[39561] = 3'b110;
        rom_memory[39562] = 3'b110;
        rom_memory[39563] = 3'b110;
        rom_memory[39564] = 3'b110;
        rom_memory[39565] = 3'b110;
        rom_memory[39566] = 3'b110;
        rom_memory[39567] = 3'b110;
        rom_memory[39568] = 3'b110;
        rom_memory[39569] = 3'b110;
        rom_memory[39570] = 3'b110;
        rom_memory[39571] = 3'b111;
        rom_memory[39572] = 3'b111;
        rom_memory[39573] = 3'b111;
        rom_memory[39574] = 3'b111;
        rom_memory[39575] = 3'b111;
        rom_memory[39576] = 3'b111;
        rom_memory[39577] = 3'b111;
        rom_memory[39578] = 3'b111;
        rom_memory[39579] = 3'b111;
        rom_memory[39580] = 3'b111;
        rom_memory[39581] = 3'b111;
        rom_memory[39582] = 3'b111;
        rom_memory[39583] = 3'b111;
        rom_memory[39584] = 3'b111;
        rom_memory[39585] = 3'b111;
        rom_memory[39586] = 3'b111;
        rom_memory[39587] = 3'b111;
        rom_memory[39588] = 3'b111;
        rom_memory[39589] = 3'b111;
        rom_memory[39590] = 3'b111;
        rom_memory[39591] = 3'b111;
        rom_memory[39592] = 3'b111;
        rom_memory[39593] = 3'b111;
        rom_memory[39594] = 3'b111;
        rom_memory[39595] = 3'b111;
        rom_memory[39596] = 3'b111;
        rom_memory[39597] = 3'b111;
        rom_memory[39598] = 3'b111;
        rom_memory[39599] = 3'b111;
        rom_memory[39600] = 3'b110;
        rom_memory[39601] = 3'b110;
        rom_memory[39602] = 3'b110;
        rom_memory[39603] = 3'b110;
        rom_memory[39604] = 3'b110;
        rom_memory[39605] = 3'b110;
        rom_memory[39606] = 3'b110;
        rom_memory[39607] = 3'b110;
        rom_memory[39608] = 3'b110;
        rom_memory[39609] = 3'b110;
        rom_memory[39610] = 3'b111;
        rom_memory[39611] = 3'b111;
        rom_memory[39612] = 3'b111;
        rom_memory[39613] = 3'b111;
        rom_memory[39614] = 3'b111;
        rom_memory[39615] = 3'b111;
        rom_memory[39616] = 3'b111;
        rom_memory[39617] = 3'b111;
        rom_memory[39618] = 3'b111;
        rom_memory[39619] = 3'b111;
        rom_memory[39620] = 3'b111;
        rom_memory[39621] = 3'b110;
        rom_memory[39622] = 3'b110;
        rom_memory[39623] = 3'b110;
        rom_memory[39624] = 3'b110;
        rom_memory[39625] = 3'b110;
        rom_memory[39626] = 3'b110;
        rom_memory[39627] = 3'b110;
        rom_memory[39628] = 3'b110;
        rom_memory[39629] = 3'b110;
        rom_memory[39630] = 3'b110;
        rom_memory[39631] = 3'b110;
        rom_memory[39632] = 3'b110;
        rom_memory[39633] = 3'b110;
        rom_memory[39634] = 3'b110;
        rom_memory[39635] = 3'b110;
        rom_memory[39636] = 3'b110;
        rom_memory[39637] = 3'b110;
        rom_memory[39638] = 3'b110;
        rom_memory[39639] = 3'b110;
        rom_memory[39640] = 3'b110;
        rom_memory[39641] = 3'b111;
        rom_memory[39642] = 3'b111;
        rom_memory[39643] = 3'b111;
        rom_memory[39644] = 3'b111;
        rom_memory[39645] = 3'b111;
        rom_memory[39646] = 3'b111;
        rom_memory[39647] = 3'b111;
        rom_memory[39648] = 3'b111;
        rom_memory[39649] = 3'b111;
        rom_memory[39650] = 3'b111;
        rom_memory[39651] = 3'b111;
        rom_memory[39652] = 3'b111;
        rom_memory[39653] = 3'b111;
        rom_memory[39654] = 3'b110;
        rom_memory[39655] = 3'b000;
        rom_memory[39656] = 3'b000;
        rom_memory[39657] = 3'b110;
        rom_memory[39658] = 3'b110;
        rom_memory[39659] = 3'b110;
        rom_memory[39660] = 3'b100;
        rom_memory[39661] = 3'b100;
        rom_memory[39662] = 3'b111;
        rom_memory[39663] = 3'b100;
        rom_memory[39664] = 3'b100;
        rom_memory[39665] = 3'b110;
        rom_memory[39666] = 3'b111;
        rom_memory[39667] = 3'b111;
        rom_memory[39668] = 3'b111;
        rom_memory[39669] = 3'b110;
        rom_memory[39670] = 3'b111;
        rom_memory[39671] = 3'b111;
        rom_memory[39672] = 3'b111;
        rom_memory[39673] = 3'b110;
        rom_memory[39674] = 3'b110;
        rom_memory[39675] = 3'b110;
        rom_memory[39676] = 3'b110;
        rom_memory[39677] = 3'b110;
        rom_memory[39678] = 3'b000;
        rom_memory[39679] = 3'b000;
        rom_memory[39680] = 3'b110;
        rom_memory[39681] = 3'b111;
        rom_memory[39682] = 3'b000;
        rom_memory[39683] = 3'b111;
        rom_memory[39684] = 3'b110;
        rom_memory[39685] = 3'b110;
        rom_memory[39686] = 3'b110;
        rom_memory[39687] = 3'b110;
        rom_memory[39688] = 3'b110;
        rom_memory[39689] = 3'b110;
        rom_memory[39690] = 3'b110;
        rom_memory[39691] = 3'b110;
        rom_memory[39692] = 3'b110;
        rom_memory[39693] = 3'b110;
        rom_memory[39694] = 3'b110;
        rom_memory[39695] = 3'b110;
        rom_memory[39696] = 3'b110;
        rom_memory[39697] = 3'b110;
        rom_memory[39698] = 3'b111;
        rom_memory[39699] = 3'b111;
        rom_memory[39700] = 3'b111;
        rom_memory[39701] = 3'b111;
        rom_memory[39702] = 3'b110;
        rom_memory[39703] = 3'b110;
        rom_memory[39704] = 3'b110;
        rom_memory[39705] = 3'b110;
        rom_memory[39706] = 3'b110;
        rom_memory[39707] = 3'b110;
        rom_memory[39708] = 3'b110;
        rom_memory[39709] = 3'b110;
        rom_memory[39710] = 3'b110;
        rom_memory[39711] = 3'b110;
        rom_memory[39712] = 3'b110;
        rom_memory[39713] = 3'b110;
        rom_memory[39714] = 3'b110;
        rom_memory[39715] = 3'b110;
        rom_memory[39716] = 3'b110;
        rom_memory[39717] = 3'b110;
        rom_memory[39718] = 3'b110;
        rom_memory[39719] = 3'b110;
        rom_memory[39720] = 3'b110;
        rom_memory[39721] = 3'b110;
        rom_memory[39722] = 3'b110;
        rom_memory[39723] = 3'b110;
        rom_memory[39724] = 3'b110;
        rom_memory[39725] = 3'b110;
        rom_memory[39726] = 3'b110;
        rom_memory[39727] = 3'b110;
        rom_memory[39728] = 3'b110;
        rom_memory[39729] = 3'b110;
        rom_memory[39730] = 3'b110;
        rom_memory[39731] = 3'b110;
        rom_memory[39732] = 3'b110;
        rom_memory[39733] = 3'b110;
        rom_memory[39734] = 3'b110;
        rom_memory[39735] = 3'b110;
        rom_memory[39736] = 3'b110;
        rom_memory[39737] = 3'b110;
        rom_memory[39738] = 3'b110;
        rom_memory[39739] = 3'b110;
        rom_memory[39740] = 3'b110;
        rom_memory[39741] = 3'b110;
        rom_memory[39742] = 3'b110;
        rom_memory[39743] = 3'b110;
        rom_memory[39744] = 3'b110;
        rom_memory[39745] = 3'b110;
        rom_memory[39746] = 3'b110;
        rom_memory[39747] = 3'b110;
        rom_memory[39748] = 3'b110;
        rom_memory[39749] = 3'b110;
        rom_memory[39750] = 3'b110;
        rom_memory[39751] = 3'b110;
        rom_memory[39752] = 3'b110;
        rom_memory[39753] = 3'b110;
        rom_memory[39754] = 3'b110;
        rom_memory[39755] = 3'b110;
        rom_memory[39756] = 3'b110;
        rom_memory[39757] = 3'b110;
        rom_memory[39758] = 3'b110;
        rom_memory[39759] = 3'b110;
        rom_memory[39760] = 3'b110;
        rom_memory[39761] = 3'b110;
        rom_memory[39762] = 3'b110;
        rom_memory[39763] = 3'b110;
        rom_memory[39764] = 3'b110;
        rom_memory[39765] = 3'b110;
        rom_memory[39766] = 3'b000;
        rom_memory[39767] = 3'b000;
        rom_memory[39768] = 3'b000;
        rom_memory[39769] = 3'b000;
        rom_memory[39770] = 3'b000;
        rom_memory[39771] = 3'b000;
        rom_memory[39772] = 3'b000;
        rom_memory[39773] = 3'b000;
        rom_memory[39774] = 3'b000;
        rom_memory[39775] = 3'b000;
        rom_memory[39776] = 3'b000;
        rom_memory[39777] = 3'b000;
        rom_memory[39778] = 3'b000;
        rom_memory[39779] = 3'b000;
        rom_memory[39780] = 3'b000;
        rom_memory[39781] = 3'b000;
        rom_memory[39782] = 3'b111;
        rom_memory[39783] = 3'b111;
        rom_memory[39784] = 3'b110;
        rom_memory[39785] = 3'b110;
        rom_memory[39786] = 3'b110;
        rom_memory[39787] = 3'b110;
        rom_memory[39788] = 3'b110;
        rom_memory[39789] = 3'b110;
        rom_memory[39790] = 3'b110;
        rom_memory[39791] = 3'b110;
        rom_memory[39792] = 3'b110;
        rom_memory[39793] = 3'b110;
        rom_memory[39794] = 3'b110;
        rom_memory[39795] = 3'b110;
        rom_memory[39796] = 3'b110;
        rom_memory[39797] = 3'b110;
        rom_memory[39798] = 3'b110;
        rom_memory[39799] = 3'b110;
        rom_memory[39800] = 3'b110;
        rom_memory[39801] = 3'b110;
        rom_memory[39802] = 3'b110;
        rom_memory[39803] = 3'b110;
        rom_memory[39804] = 3'b110;
        rom_memory[39805] = 3'b110;
        rom_memory[39806] = 3'b110;
        rom_memory[39807] = 3'b110;
        rom_memory[39808] = 3'b110;
        rom_memory[39809] = 3'b110;
        rom_memory[39810] = 3'b110;
        rom_memory[39811] = 3'b110;
        rom_memory[39812] = 3'b110;
        rom_memory[39813] = 3'b111;
        rom_memory[39814] = 3'b111;
        rom_memory[39815] = 3'b111;
        rom_memory[39816] = 3'b111;
        rom_memory[39817] = 3'b111;
        rom_memory[39818] = 3'b111;
        rom_memory[39819] = 3'b111;
        rom_memory[39820] = 3'b111;
        rom_memory[39821] = 3'b111;
        rom_memory[39822] = 3'b111;
        rom_memory[39823] = 3'b111;
        rom_memory[39824] = 3'b111;
        rom_memory[39825] = 3'b111;
        rom_memory[39826] = 3'b111;
        rom_memory[39827] = 3'b111;
        rom_memory[39828] = 3'b111;
        rom_memory[39829] = 3'b111;
        rom_memory[39830] = 3'b111;
        rom_memory[39831] = 3'b111;
        rom_memory[39832] = 3'b111;
        rom_memory[39833] = 3'b111;
        rom_memory[39834] = 3'b111;
        rom_memory[39835] = 3'b111;
        rom_memory[39836] = 3'b111;
        rom_memory[39837] = 3'b111;
        rom_memory[39838] = 3'b111;
        rom_memory[39839] = 3'b111;
        rom_memory[39840] = 3'b110;
        rom_memory[39841] = 3'b110;
        rom_memory[39842] = 3'b110;
        rom_memory[39843] = 3'b110;
        rom_memory[39844] = 3'b110;
        rom_memory[39845] = 3'b110;
        rom_memory[39846] = 3'b110;
        rom_memory[39847] = 3'b110;
        rom_memory[39848] = 3'b110;
        rom_memory[39849] = 3'b110;
        rom_memory[39850] = 3'b111;
        rom_memory[39851] = 3'b111;
        rom_memory[39852] = 3'b111;
        rom_memory[39853] = 3'b111;
        rom_memory[39854] = 3'b111;
        rom_memory[39855] = 3'b111;
        rom_memory[39856] = 3'b111;
        rom_memory[39857] = 3'b111;
        rom_memory[39858] = 3'b111;
        rom_memory[39859] = 3'b111;
        rom_memory[39860] = 3'b111;
        rom_memory[39861] = 3'b110;
        rom_memory[39862] = 3'b110;
        rom_memory[39863] = 3'b110;
        rom_memory[39864] = 3'b110;
        rom_memory[39865] = 3'b110;
        rom_memory[39866] = 3'b110;
        rom_memory[39867] = 3'b110;
        rom_memory[39868] = 3'b110;
        rom_memory[39869] = 3'b110;
        rom_memory[39870] = 3'b110;
        rom_memory[39871] = 3'b110;
        rom_memory[39872] = 3'b110;
        rom_memory[39873] = 3'b110;
        rom_memory[39874] = 3'b110;
        rom_memory[39875] = 3'b110;
        rom_memory[39876] = 3'b110;
        rom_memory[39877] = 3'b110;
        rom_memory[39878] = 3'b110;
        rom_memory[39879] = 3'b110;
        rom_memory[39880] = 3'b110;
        rom_memory[39881] = 3'b111;
        rom_memory[39882] = 3'b111;
        rom_memory[39883] = 3'b111;
        rom_memory[39884] = 3'b111;
        rom_memory[39885] = 3'b111;
        rom_memory[39886] = 3'b111;
        rom_memory[39887] = 3'b111;
        rom_memory[39888] = 3'b111;
        rom_memory[39889] = 3'b111;
        rom_memory[39890] = 3'b111;
        rom_memory[39891] = 3'b111;
        rom_memory[39892] = 3'b111;
        rom_memory[39893] = 3'b111;
        rom_memory[39894] = 3'b010;
        rom_memory[39895] = 3'b000;
        rom_memory[39896] = 3'b010;
        rom_memory[39897] = 3'b111;
        rom_memory[39898] = 3'b111;
        rom_memory[39899] = 3'b000;
        rom_memory[39900] = 3'b000;
        rom_memory[39901] = 3'b100;
        rom_memory[39902] = 3'b111;
        rom_memory[39903] = 3'b000;
        rom_memory[39904] = 3'b000;
        rom_memory[39905] = 3'b000;
        rom_memory[39906] = 3'b100;
        rom_memory[39907] = 3'b100;
        rom_memory[39908] = 3'b110;
        rom_memory[39909] = 3'b111;
        rom_memory[39910] = 3'b110;
        rom_memory[39911] = 3'b110;
        rom_memory[39912] = 3'b111;
        rom_memory[39913] = 3'b110;
        rom_memory[39914] = 3'b111;
        rom_memory[39915] = 3'b111;
        rom_memory[39916] = 3'b111;
        rom_memory[39917] = 3'b100;
        rom_memory[39918] = 3'b000;
        rom_memory[39919] = 3'b110;
        rom_memory[39920] = 3'b100;
        rom_memory[39921] = 3'b000;
        rom_memory[39922] = 3'b100;
        rom_memory[39923] = 3'b110;
        rom_memory[39924] = 3'b110;
        rom_memory[39925] = 3'b110;
        rom_memory[39926] = 3'b110;
        rom_memory[39927] = 3'b110;
        rom_memory[39928] = 3'b110;
        rom_memory[39929] = 3'b110;
        rom_memory[39930] = 3'b110;
        rom_memory[39931] = 3'b110;
        rom_memory[39932] = 3'b110;
        rom_memory[39933] = 3'b110;
        rom_memory[39934] = 3'b110;
        rom_memory[39935] = 3'b110;
        rom_memory[39936] = 3'b110;
        rom_memory[39937] = 3'b110;
        rom_memory[39938] = 3'b110;
        rom_memory[39939] = 3'b110;
        rom_memory[39940] = 3'b110;
        rom_memory[39941] = 3'b110;
        rom_memory[39942] = 3'b110;
        rom_memory[39943] = 3'b110;
        rom_memory[39944] = 3'b110;
        rom_memory[39945] = 3'b110;
        rom_memory[39946] = 3'b110;
        rom_memory[39947] = 3'b110;
        rom_memory[39948] = 3'b110;
        rom_memory[39949] = 3'b110;
        rom_memory[39950] = 3'b110;
        rom_memory[39951] = 3'b110;
        rom_memory[39952] = 3'b110;
        rom_memory[39953] = 3'b110;
        rom_memory[39954] = 3'b110;
        rom_memory[39955] = 3'b110;
        rom_memory[39956] = 3'b110;
        rom_memory[39957] = 3'b110;
        rom_memory[39958] = 3'b110;
        rom_memory[39959] = 3'b110;
        rom_memory[39960] = 3'b110;
        rom_memory[39961] = 3'b110;
        rom_memory[39962] = 3'b110;
        rom_memory[39963] = 3'b110;
        rom_memory[39964] = 3'b110;
        rom_memory[39965] = 3'b110;
        rom_memory[39966] = 3'b110;
        rom_memory[39967] = 3'b110;
        rom_memory[39968] = 3'b110;
        rom_memory[39969] = 3'b110;
        rom_memory[39970] = 3'b110;
        rom_memory[39971] = 3'b110;
        rom_memory[39972] = 3'b110;
        rom_memory[39973] = 3'b110;
        rom_memory[39974] = 3'b110;
        rom_memory[39975] = 3'b110;
        rom_memory[39976] = 3'b110;
        rom_memory[39977] = 3'b110;
        rom_memory[39978] = 3'b110;
        rom_memory[39979] = 3'b110;
        rom_memory[39980] = 3'b110;
        rom_memory[39981] = 3'b110;
        rom_memory[39982] = 3'b110;
        rom_memory[39983] = 3'b110;
        rom_memory[39984] = 3'b110;
        rom_memory[39985] = 3'b110;
        rom_memory[39986] = 3'b110;
        rom_memory[39987] = 3'b110;
        rom_memory[39988] = 3'b110;
        rom_memory[39989] = 3'b110;
        rom_memory[39990] = 3'b110;
        rom_memory[39991] = 3'b110;
        rom_memory[39992] = 3'b110;
        rom_memory[39993] = 3'b110;
        rom_memory[39994] = 3'b110;
        rom_memory[39995] = 3'b110;
        rom_memory[39996] = 3'b110;
        rom_memory[39997] = 3'b110;
        rom_memory[39998] = 3'b110;
        rom_memory[39999] = 3'b110;
        rom_memory[40000] = 3'b110;
        rom_memory[40001] = 3'b110;
        rom_memory[40002] = 3'b110;
        rom_memory[40003] = 3'b110;
        rom_memory[40004] = 3'b110;
        rom_memory[40005] = 3'b110;
        rom_memory[40006] = 3'b110;
        rom_memory[40007] = 3'b100;
        rom_memory[40008] = 3'b000;
        rom_memory[40009] = 3'b000;
        rom_memory[40010] = 3'b000;
        rom_memory[40011] = 3'b000;
        rom_memory[40012] = 3'b000;
        rom_memory[40013] = 3'b000;
        rom_memory[40014] = 3'b000;
        rom_memory[40015] = 3'b000;
        rom_memory[40016] = 3'b000;
        rom_memory[40017] = 3'b000;
        rom_memory[40018] = 3'b000;
        rom_memory[40019] = 3'b000;
        rom_memory[40020] = 3'b000;
        rom_memory[40021] = 3'b000;
        rom_memory[40022] = 3'b000;
        rom_memory[40023] = 3'b110;
        rom_memory[40024] = 3'b111;
        rom_memory[40025] = 3'b111;
        rom_memory[40026] = 3'b110;
        rom_memory[40027] = 3'b110;
        rom_memory[40028] = 3'b110;
        rom_memory[40029] = 3'b110;
        rom_memory[40030] = 3'b110;
        rom_memory[40031] = 3'b110;
        rom_memory[40032] = 3'b110;
        rom_memory[40033] = 3'b110;
        rom_memory[40034] = 3'b110;
        rom_memory[40035] = 3'b110;
        rom_memory[40036] = 3'b110;
        rom_memory[40037] = 3'b110;
        rom_memory[40038] = 3'b110;
        rom_memory[40039] = 3'b110;
        rom_memory[40040] = 3'b110;
        rom_memory[40041] = 3'b110;
        rom_memory[40042] = 3'b110;
        rom_memory[40043] = 3'b110;
        rom_memory[40044] = 3'b110;
        rom_memory[40045] = 3'b110;
        rom_memory[40046] = 3'b110;
        rom_memory[40047] = 3'b110;
        rom_memory[40048] = 3'b110;
        rom_memory[40049] = 3'b110;
        rom_memory[40050] = 3'b110;
        rom_memory[40051] = 3'b110;
        rom_memory[40052] = 3'b110;
        rom_memory[40053] = 3'b110;
        rom_memory[40054] = 3'b110;
        rom_memory[40055] = 3'b111;
        rom_memory[40056] = 3'b110;
        rom_memory[40057] = 3'b111;
        rom_memory[40058] = 3'b111;
        rom_memory[40059] = 3'b111;
        rom_memory[40060] = 3'b111;
        rom_memory[40061] = 3'b111;
        rom_memory[40062] = 3'b111;
        rom_memory[40063] = 3'b111;
        rom_memory[40064] = 3'b111;
        rom_memory[40065] = 3'b111;
        rom_memory[40066] = 3'b111;
        rom_memory[40067] = 3'b111;
        rom_memory[40068] = 3'b111;
        rom_memory[40069] = 3'b111;
        rom_memory[40070] = 3'b111;
        rom_memory[40071] = 3'b111;
        rom_memory[40072] = 3'b111;
        rom_memory[40073] = 3'b111;
        rom_memory[40074] = 3'b111;
        rom_memory[40075] = 3'b111;
        rom_memory[40076] = 3'b111;
        rom_memory[40077] = 3'b111;
        rom_memory[40078] = 3'b111;
        rom_memory[40079] = 3'b111;
        rom_memory[40080] = 3'b110;
        rom_memory[40081] = 3'b110;
        rom_memory[40082] = 3'b110;
        rom_memory[40083] = 3'b110;
        rom_memory[40084] = 3'b110;
        rom_memory[40085] = 3'b110;
        rom_memory[40086] = 3'b110;
        rom_memory[40087] = 3'b110;
        rom_memory[40088] = 3'b110;
        rom_memory[40089] = 3'b110;
        rom_memory[40090] = 3'b110;
        rom_memory[40091] = 3'b111;
        rom_memory[40092] = 3'b111;
        rom_memory[40093] = 3'b111;
        rom_memory[40094] = 3'b111;
        rom_memory[40095] = 3'b111;
        rom_memory[40096] = 3'b111;
        rom_memory[40097] = 3'b111;
        rom_memory[40098] = 3'b111;
        rom_memory[40099] = 3'b111;
        rom_memory[40100] = 3'b111;
        rom_memory[40101] = 3'b110;
        rom_memory[40102] = 3'b110;
        rom_memory[40103] = 3'b110;
        rom_memory[40104] = 3'b110;
        rom_memory[40105] = 3'b110;
        rom_memory[40106] = 3'b110;
        rom_memory[40107] = 3'b110;
        rom_memory[40108] = 3'b110;
        rom_memory[40109] = 3'b110;
        rom_memory[40110] = 3'b110;
        rom_memory[40111] = 3'b110;
        rom_memory[40112] = 3'b110;
        rom_memory[40113] = 3'b110;
        rom_memory[40114] = 3'b110;
        rom_memory[40115] = 3'b110;
        rom_memory[40116] = 3'b110;
        rom_memory[40117] = 3'b110;
        rom_memory[40118] = 3'b110;
        rom_memory[40119] = 3'b111;
        rom_memory[40120] = 3'b111;
        rom_memory[40121] = 3'b111;
        rom_memory[40122] = 3'b111;
        rom_memory[40123] = 3'b111;
        rom_memory[40124] = 3'b111;
        rom_memory[40125] = 3'b111;
        rom_memory[40126] = 3'b111;
        rom_memory[40127] = 3'b111;
        rom_memory[40128] = 3'b111;
        rom_memory[40129] = 3'b111;
        rom_memory[40130] = 3'b111;
        rom_memory[40131] = 3'b111;
        rom_memory[40132] = 3'b111;
        rom_memory[40133] = 3'b110;
        rom_memory[40134] = 3'b010;
        rom_memory[40135] = 3'b000;
        rom_memory[40136] = 3'b110;
        rom_memory[40137] = 3'b111;
        rom_memory[40138] = 3'b111;
        rom_memory[40139] = 3'b000;
        rom_memory[40140] = 3'b000;
        rom_memory[40141] = 3'b110;
        rom_memory[40142] = 3'b110;
        rom_memory[40143] = 3'b110;
        rom_memory[40144] = 3'b100;
        rom_memory[40145] = 3'b000;
        rom_memory[40146] = 3'b000;
        rom_memory[40147] = 3'b100;
        rom_memory[40148] = 3'b111;
        rom_memory[40149] = 3'b111;
        rom_memory[40150] = 3'b110;
        rom_memory[40151] = 3'b100;
        rom_memory[40152] = 3'b111;
        rom_memory[40153] = 3'b111;
        rom_memory[40154] = 3'b111;
        rom_memory[40155] = 3'b111;
        rom_memory[40156] = 3'b111;
        rom_memory[40157] = 3'b110;
        rom_memory[40158] = 3'b000;
        rom_memory[40159] = 3'b111;
        rom_memory[40160] = 3'b000;
        rom_memory[40161] = 3'b000;
        rom_memory[40162] = 3'b100;
        rom_memory[40163] = 3'b110;
        rom_memory[40164] = 3'b110;
        rom_memory[40165] = 3'b110;
        rom_memory[40166] = 3'b110;
        rom_memory[40167] = 3'b110;
        rom_memory[40168] = 3'b110;
        rom_memory[40169] = 3'b110;
        rom_memory[40170] = 3'b110;
        rom_memory[40171] = 3'b110;
        rom_memory[40172] = 3'b110;
        rom_memory[40173] = 3'b110;
        rom_memory[40174] = 3'b110;
        rom_memory[40175] = 3'b110;
        rom_memory[40176] = 3'b110;
        rom_memory[40177] = 3'b110;
        rom_memory[40178] = 3'b110;
        rom_memory[40179] = 3'b110;
        rom_memory[40180] = 3'b110;
        rom_memory[40181] = 3'b110;
        rom_memory[40182] = 3'b110;
        rom_memory[40183] = 3'b110;
        rom_memory[40184] = 3'b110;
        rom_memory[40185] = 3'b110;
        rom_memory[40186] = 3'b110;
        rom_memory[40187] = 3'b110;
        rom_memory[40188] = 3'b110;
        rom_memory[40189] = 3'b110;
        rom_memory[40190] = 3'b110;
        rom_memory[40191] = 3'b110;
        rom_memory[40192] = 3'b110;
        rom_memory[40193] = 3'b110;
        rom_memory[40194] = 3'b110;
        rom_memory[40195] = 3'b110;
        rom_memory[40196] = 3'b110;
        rom_memory[40197] = 3'b110;
        rom_memory[40198] = 3'b110;
        rom_memory[40199] = 3'b110;
        rom_memory[40200] = 3'b110;
        rom_memory[40201] = 3'b110;
        rom_memory[40202] = 3'b110;
        rom_memory[40203] = 3'b110;
        rom_memory[40204] = 3'b110;
        rom_memory[40205] = 3'b110;
        rom_memory[40206] = 3'b110;
        rom_memory[40207] = 3'b110;
        rom_memory[40208] = 3'b110;
        rom_memory[40209] = 3'b110;
        rom_memory[40210] = 3'b110;
        rom_memory[40211] = 3'b110;
        rom_memory[40212] = 3'b110;
        rom_memory[40213] = 3'b110;
        rom_memory[40214] = 3'b110;
        rom_memory[40215] = 3'b110;
        rom_memory[40216] = 3'b110;
        rom_memory[40217] = 3'b110;
        rom_memory[40218] = 3'b110;
        rom_memory[40219] = 3'b110;
        rom_memory[40220] = 3'b110;
        rom_memory[40221] = 3'b110;
        rom_memory[40222] = 3'b110;
        rom_memory[40223] = 3'b110;
        rom_memory[40224] = 3'b110;
        rom_memory[40225] = 3'b110;
        rom_memory[40226] = 3'b110;
        rom_memory[40227] = 3'b110;
        rom_memory[40228] = 3'b110;
        rom_memory[40229] = 3'b110;
        rom_memory[40230] = 3'b110;
        rom_memory[40231] = 3'b110;
        rom_memory[40232] = 3'b110;
        rom_memory[40233] = 3'b110;
        rom_memory[40234] = 3'b110;
        rom_memory[40235] = 3'b110;
        rom_memory[40236] = 3'b110;
        rom_memory[40237] = 3'b110;
        rom_memory[40238] = 3'b110;
        rom_memory[40239] = 3'b110;
        rom_memory[40240] = 3'b110;
        rom_memory[40241] = 3'b110;
        rom_memory[40242] = 3'b110;
        rom_memory[40243] = 3'b110;
        rom_memory[40244] = 3'b110;
        rom_memory[40245] = 3'b110;
        rom_memory[40246] = 3'b110;
        rom_memory[40247] = 3'b110;
        rom_memory[40248] = 3'b110;
        rom_memory[40249] = 3'b000;
        rom_memory[40250] = 3'b000;
        rom_memory[40251] = 3'b000;
        rom_memory[40252] = 3'b000;
        rom_memory[40253] = 3'b000;
        rom_memory[40254] = 3'b000;
        rom_memory[40255] = 3'b000;
        rom_memory[40256] = 3'b000;
        rom_memory[40257] = 3'b000;
        rom_memory[40258] = 3'b000;
        rom_memory[40259] = 3'b000;
        rom_memory[40260] = 3'b000;
        rom_memory[40261] = 3'b000;
        rom_memory[40262] = 3'b000;
        rom_memory[40263] = 3'b000;
        rom_memory[40264] = 3'b100;
        rom_memory[40265] = 3'b111;
        rom_memory[40266] = 3'b111;
        rom_memory[40267] = 3'b110;
        rom_memory[40268] = 3'b110;
        rom_memory[40269] = 3'b110;
        rom_memory[40270] = 3'b110;
        rom_memory[40271] = 3'b110;
        rom_memory[40272] = 3'b110;
        rom_memory[40273] = 3'b110;
        rom_memory[40274] = 3'b110;
        rom_memory[40275] = 3'b110;
        rom_memory[40276] = 3'b110;
        rom_memory[40277] = 3'b110;
        rom_memory[40278] = 3'b110;
        rom_memory[40279] = 3'b110;
        rom_memory[40280] = 3'b110;
        rom_memory[40281] = 3'b110;
        rom_memory[40282] = 3'b110;
        rom_memory[40283] = 3'b110;
        rom_memory[40284] = 3'b110;
        rom_memory[40285] = 3'b110;
        rom_memory[40286] = 3'b110;
        rom_memory[40287] = 3'b110;
        rom_memory[40288] = 3'b110;
        rom_memory[40289] = 3'b110;
        rom_memory[40290] = 3'b110;
        rom_memory[40291] = 3'b110;
        rom_memory[40292] = 3'b110;
        rom_memory[40293] = 3'b110;
        rom_memory[40294] = 3'b110;
        rom_memory[40295] = 3'b111;
        rom_memory[40296] = 3'b110;
        rom_memory[40297] = 3'b111;
        rom_memory[40298] = 3'b111;
        rom_memory[40299] = 3'b111;
        rom_memory[40300] = 3'b111;
        rom_memory[40301] = 3'b111;
        rom_memory[40302] = 3'b111;
        rom_memory[40303] = 3'b111;
        rom_memory[40304] = 3'b111;
        rom_memory[40305] = 3'b111;
        rom_memory[40306] = 3'b111;
        rom_memory[40307] = 3'b111;
        rom_memory[40308] = 3'b111;
        rom_memory[40309] = 3'b111;
        rom_memory[40310] = 3'b111;
        rom_memory[40311] = 3'b111;
        rom_memory[40312] = 3'b111;
        rom_memory[40313] = 3'b111;
        rom_memory[40314] = 3'b111;
        rom_memory[40315] = 3'b111;
        rom_memory[40316] = 3'b111;
        rom_memory[40317] = 3'b111;
        rom_memory[40318] = 3'b111;
        rom_memory[40319] = 3'b111;
        rom_memory[40320] = 3'b110;
        rom_memory[40321] = 3'b110;
        rom_memory[40322] = 3'b110;
        rom_memory[40323] = 3'b110;
        rom_memory[40324] = 3'b110;
        rom_memory[40325] = 3'b110;
        rom_memory[40326] = 3'b110;
        rom_memory[40327] = 3'b110;
        rom_memory[40328] = 3'b110;
        rom_memory[40329] = 3'b110;
        rom_memory[40330] = 3'b111;
        rom_memory[40331] = 3'b111;
        rom_memory[40332] = 3'b111;
        rom_memory[40333] = 3'b111;
        rom_memory[40334] = 3'b111;
        rom_memory[40335] = 3'b111;
        rom_memory[40336] = 3'b111;
        rom_memory[40337] = 3'b111;
        rom_memory[40338] = 3'b111;
        rom_memory[40339] = 3'b111;
        rom_memory[40340] = 3'b111;
        rom_memory[40341] = 3'b110;
        rom_memory[40342] = 3'b110;
        rom_memory[40343] = 3'b110;
        rom_memory[40344] = 3'b110;
        rom_memory[40345] = 3'b110;
        rom_memory[40346] = 3'b110;
        rom_memory[40347] = 3'b110;
        rom_memory[40348] = 3'b110;
        rom_memory[40349] = 3'b110;
        rom_memory[40350] = 3'b110;
        rom_memory[40351] = 3'b110;
        rom_memory[40352] = 3'b110;
        rom_memory[40353] = 3'b110;
        rom_memory[40354] = 3'b110;
        rom_memory[40355] = 3'b110;
        rom_memory[40356] = 3'b110;
        rom_memory[40357] = 3'b110;
        rom_memory[40358] = 3'b110;
        rom_memory[40359] = 3'b111;
        rom_memory[40360] = 3'b111;
        rom_memory[40361] = 3'b111;
        rom_memory[40362] = 3'b111;
        rom_memory[40363] = 3'b111;
        rom_memory[40364] = 3'b111;
        rom_memory[40365] = 3'b111;
        rom_memory[40366] = 3'b111;
        rom_memory[40367] = 3'b111;
        rom_memory[40368] = 3'b111;
        rom_memory[40369] = 3'b111;
        rom_memory[40370] = 3'b111;
        rom_memory[40371] = 3'b111;
        rom_memory[40372] = 3'b111;
        rom_memory[40373] = 3'b110;
        rom_memory[40374] = 3'b010;
        rom_memory[40375] = 3'b010;
        rom_memory[40376] = 3'b110;
        rom_memory[40377] = 3'b111;
        rom_memory[40378] = 3'b111;
        rom_memory[40379] = 3'b000;
        rom_memory[40380] = 3'b000;
        rom_memory[40381] = 3'b100;
        rom_memory[40382] = 3'b110;
        rom_memory[40383] = 3'b110;
        rom_memory[40384] = 3'b110;
        rom_memory[40385] = 3'b110;
        rom_memory[40386] = 3'b100;
        rom_memory[40387] = 3'b000;
        rom_memory[40388] = 3'b100;
        rom_memory[40389] = 3'b100;
        rom_memory[40390] = 3'b100;
        rom_memory[40391] = 3'b111;
        rom_memory[40392] = 3'b111;
        rom_memory[40393] = 3'b111;
        rom_memory[40394] = 3'b110;
        rom_memory[40395] = 3'b110;
        rom_memory[40396] = 3'b110;
        rom_memory[40397] = 3'b100;
        rom_memory[40398] = 3'b000;
        rom_memory[40399] = 3'b110;
        rom_memory[40400] = 3'b100;
        rom_memory[40401] = 3'b000;
        rom_memory[40402] = 3'b110;
        rom_memory[40403] = 3'b110;
        rom_memory[40404] = 3'b110;
        rom_memory[40405] = 3'b110;
        rom_memory[40406] = 3'b110;
        rom_memory[40407] = 3'b110;
        rom_memory[40408] = 3'b110;
        rom_memory[40409] = 3'b110;
        rom_memory[40410] = 3'b110;
        rom_memory[40411] = 3'b110;
        rom_memory[40412] = 3'b110;
        rom_memory[40413] = 3'b110;
        rom_memory[40414] = 3'b110;
        rom_memory[40415] = 3'b110;
        rom_memory[40416] = 3'b110;
        rom_memory[40417] = 3'b110;
        rom_memory[40418] = 3'b110;
        rom_memory[40419] = 3'b110;
        rom_memory[40420] = 3'b110;
        rom_memory[40421] = 3'b110;
        rom_memory[40422] = 3'b111;
        rom_memory[40423] = 3'b111;
        rom_memory[40424] = 3'b111;
        rom_memory[40425] = 3'b111;
        rom_memory[40426] = 3'b110;
        rom_memory[40427] = 3'b110;
        rom_memory[40428] = 3'b110;
        rom_memory[40429] = 3'b110;
        rom_memory[40430] = 3'b110;
        rom_memory[40431] = 3'b110;
        rom_memory[40432] = 3'b110;
        rom_memory[40433] = 3'b110;
        rom_memory[40434] = 3'b110;
        rom_memory[40435] = 3'b110;
        rom_memory[40436] = 3'b110;
        rom_memory[40437] = 3'b110;
        rom_memory[40438] = 3'b110;
        rom_memory[40439] = 3'b110;
        rom_memory[40440] = 3'b110;
        rom_memory[40441] = 3'b110;
        rom_memory[40442] = 3'b110;
        rom_memory[40443] = 3'b110;
        rom_memory[40444] = 3'b110;
        rom_memory[40445] = 3'b110;
        rom_memory[40446] = 3'b110;
        rom_memory[40447] = 3'b110;
        rom_memory[40448] = 3'b110;
        rom_memory[40449] = 3'b110;
        rom_memory[40450] = 3'b110;
        rom_memory[40451] = 3'b110;
        rom_memory[40452] = 3'b110;
        rom_memory[40453] = 3'b110;
        rom_memory[40454] = 3'b110;
        rom_memory[40455] = 3'b110;
        rom_memory[40456] = 3'b110;
        rom_memory[40457] = 3'b110;
        rom_memory[40458] = 3'b110;
        rom_memory[40459] = 3'b110;
        rom_memory[40460] = 3'b110;
        rom_memory[40461] = 3'b110;
        rom_memory[40462] = 3'b110;
        rom_memory[40463] = 3'b110;
        rom_memory[40464] = 3'b110;
        rom_memory[40465] = 3'b110;
        rom_memory[40466] = 3'b110;
        rom_memory[40467] = 3'b110;
        rom_memory[40468] = 3'b110;
        rom_memory[40469] = 3'b110;
        rom_memory[40470] = 3'b110;
        rom_memory[40471] = 3'b110;
        rom_memory[40472] = 3'b110;
        rom_memory[40473] = 3'b110;
        rom_memory[40474] = 3'b110;
        rom_memory[40475] = 3'b110;
        rom_memory[40476] = 3'b110;
        rom_memory[40477] = 3'b110;
        rom_memory[40478] = 3'b110;
        rom_memory[40479] = 3'b110;
        rom_memory[40480] = 3'b110;
        rom_memory[40481] = 3'b110;
        rom_memory[40482] = 3'b110;
        rom_memory[40483] = 3'b110;
        rom_memory[40484] = 3'b110;
        rom_memory[40485] = 3'b110;
        rom_memory[40486] = 3'b110;
        rom_memory[40487] = 3'b110;
        rom_memory[40488] = 3'b110;
        rom_memory[40489] = 3'b110;
        rom_memory[40490] = 3'b110;
        rom_memory[40491] = 3'b000;
        rom_memory[40492] = 3'b000;
        rom_memory[40493] = 3'b000;
        rom_memory[40494] = 3'b000;
        rom_memory[40495] = 3'b000;
        rom_memory[40496] = 3'b000;
        rom_memory[40497] = 3'b000;
        rom_memory[40498] = 3'b000;
        rom_memory[40499] = 3'b000;
        rom_memory[40500] = 3'b000;
        rom_memory[40501] = 3'b000;
        rom_memory[40502] = 3'b000;
        rom_memory[40503] = 3'b000;
        rom_memory[40504] = 3'b000;
        rom_memory[40505] = 3'b000;
        rom_memory[40506] = 3'b111;
        rom_memory[40507] = 3'b111;
        rom_memory[40508] = 3'b110;
        rom_memory[40509] = 3'b110;
        rom_memory[40510] = 3'b110;
        rom_memory[40511] = 3'b110;
        rom_memory[40512] = 3'b110;
        rom_memory[40513] = 3'b110;
        rom_memory[40514] = 3'b110;
        rom_memory[40515] = 3'b110;
        rom_memory[40516] = 3'b110;
        rom_memory[40517] = 3'b110;
        rom_memory[40518] = 3'b110;
        rom_memory[40519] = 3'b110;
        rom_memory[40520] = 3'b110;
        rom_memory[40521] = 3'b110;
        rom_memory[40522] = 3'b110;
        rom_memory[40523] = 3'b110;
        rom_memory[40524] = 3'b110;
        rom_memory[40525] = 3'b110;
        rom_memory[40526] = 3'b110;
        rom_memory[40527] = 3'b110;
        rom_memory[40528] = 3'b110;
        rom_memory[40529] = 3'b110;
        rom_memory[40530] = 3'b110;
        rom_memory[40531] = 3'b110;
        rom_memory[40532] = 3'b110;
        rom_memory[40533] = 3'b110;
        rom_memory[40534] = 3'b110;
        rom_memory[40535] = 3'b110;
        rom_memory[40536] = 3'b110;
        rom_memory[40537] = 3'b110;
        rom_memory[40538] = 3'b111;
        rom_memory[40539] = 3'b111;
        rom_memory[40540] = 3'b111;
        rom_memory[40541] = 3'b111;
        rom_memory[40542] = 3'b110;
        rom_memory[40543] = 3'b111;
        rom_memory[40544] = 3'b111;
        rom_memory[40545] = 3'b111;
        rom_memory[40546] = 3'b111;
        rom_memory[40547] = 3'b111;
        rom_memory[40548] = 3'b111;
        rom_memory[40549] = 3'b111;
        rom_memory[40550] = 3'b111;
        rom_memory[40551] = 3'b111;
        rom_memory[40552] = 3'b111;
        rom_memory[40553] = 3'b111;
        rom_memory[40554] = 3'b111;
        rom_memory[40555] = 3'b111;
        rom_memory[40556] = 3'b111;
        rom_memory[40557] = 3'b111;
        rom_memory[40558] = 3'b111;
        rom_memory[40559] = 3'b111;
        rom_memory[40560] = 3'b110;
        rom_memory[40561] = 3'b110;
        rom_memory[40562] = 3'b110;
        rom_memory[40563] = 3'b110;
        rom_memory[40564] = 3'b110;
        rom_memory[40565] = 3'b110;
        rom_memory[40566] = 3'b110;
        rom_memory[40567] = 3'b110;
        rom_memory[40568] = 3'b110;
        rom_memory[40569] = 3'b110;
        rom_memory[40570] = 3'b111;
        rom_memory[40571] = 3'b111;
        rom_memory[40572] = 3'b111;
        rom_memory[40573] = 3'b111;
        rom_memory[40574] = 3'b111;
        rom_memory[40575] = 3'b111;
        rom_memory[40576] = 3'b111;
        rom_memory[40577] = 3'b111;
        rom_memory[40578] = 3'b111;
        rom_memory[40579] = 3'b111;
        rom_memory[40580] = 3'b111;
        rom_memory[40581] = 3'b110;
        rom_memory[40582] = 3'b110;
        rom_memory[40583] = 3'b110;
        rom_memory[40584] = 3'b110;
        rom_memory[40585] = 3'b110;
        rom_memory[40586] = 3'b110;
        rom_memory[40587] = 3'b110;
        rom_memory[40588] = 3'b110;
        rom_memory[40589] = 3'b110;
        rom_memory[40590] = 3'b110;
        rom_memory[40591] = 3'b110;
        rom_memory[40592] = 3'b110;
        rom_memory[40593] = 3'b110;
        rom_memory[40594] = 3'b110;
        rom_memory[40595] = 3'b110;
        rom_memory[40596] = 3'b110;
        rom_memory[40597] = 3'b110;
        rom_memory[40598] = 3'b110;
        rom_memory[40599] = 3'b111;
        rom_memory[40600] = 3'b111;
        rom_memory[40601] = 3'b111;
        rom_memory[40602] = 3'b111;
        rom_memory[40603] = 3'b111;
        rom_memory[40604] = 3'b111;
        rom_memory[40605] = 3'b111;
        rom_memory[40606] = 3'b111;
        rom_memory[40607] = 3'b111;
        rom_memory[40608] = 3'b111;
        rom_memory[40609] = 3'b111;
        rom_memory[40610] = 3'b111;
        rom_memory[40611] = 3'b111;
        rom_memory[40612] = 3'b111;
        rom_memory[40613] = 3'b110;
        rom_memory[40614] = 3'b010;
        rom_memory[40615] = 3'b110;
        rom_memory[40616] = 3'b110;
        rom_memory[40617] = 3'b111;
        rom_memory[40618] = 3'b111;
        rom_memory[40619] = 3'b000;
        rom_memory[40620] = 3'b000;
        rom_memory[40621] = 3'b010;
        rom_memory[40622] = 3'b110;
        rom_memory[40623] = 3'b110;
        rom_memory[40624] = 3'b110;
        rom_memory[40625] = 3'b110;
        rom_memory[40626] = 3'b110;
        rom_memory[40627] = 3'b100;
        rom_memory[40628] = 3'b110;
        rom_memory[40629] = 3'b000;
        rom_memory[40630] = 3'b100;
        rom_memory[40631] = 3'b111;
        rom_memory[40632] = 3'b111;
        rom_memory[40633] = 3'b111;
        rom_memory[40634] = 3'b100;
        rom_memory[40635] = 3'b100;
        rom_memory[40636] = 3'b111;
        rom_memory[40637] = 3'b111;
        rom_memory[40638] = 3'b100;
        rom_memory[40639] = 3'b000;
        rom_memory[40640] = 3'b100;
        rom_memory[40641] = 3'b110;
        rom_memory[40642] = 3'b110;
        rom_memory[40643] = 3'b110;
        rom_memory[40644] = 3'b110;
        rom_memory[40645] = 3'b110;
        rom_memory[40646] = 3'b110;
        rom_memory[40647] = 3'b111;
        rom_memory[40648] = 3'b110;
        rom_memory[40649] = 3'b110;
        rom_memory[40650] = 3'b111;
        rom_memory[40651] = 3'b111;
        rom_memory[40652] = 3'b110;
        rom_memory[40653] = 3'b110;
        rom_memory[40654] = 3'b110;
        rom_memory[40655] = 3'b110;
        rom_memory[40656] = 3'b110;
        rom_memory[40657] = 3'b110;
        rom_memory[40658] = 3'b110;
        rom_memory[40659] = 3'b110;
        rom_memory[40660] = 3'b110;
        rom_memory[40661] = 3'b110;
        rom_memory[40662] = 3'b111;
        rom_memory[40663] = 3'b111;
        rom_memory[40664] = 3'b111;
        rom_memory[40665] = 3'b111;
        rom_memory[40666] = 3'b111;
        rom_memory[40667] = 3'b110;
        rom_memory[40668] = 3'b110;
        rom_memory[40669] = 3'b110;
        rom_memory[40670] = 3'b110;
        rom_memory[40671] = 3'b110;
        rom_memory[40672] = 3'b110;
        rom_memory[40673] = 3'b110;
        rom_memory[40674] = 3'b110;
        rom_memory[40675] = 3'b110;
        rom_memory[40676] = 3'b110;
        rom_memory[40677] = 3'b110;
        rom_memory[40678] = 3'b110;
        rom_memory[40679] = 3'b110;
        rom_memory[40680] = 3'b110;
        rom_memory[40681] = 3'b110;
        rom_memory[40682] = 3'b110;
        rom_memory[40683] = 3'b110;
        rom_memory[40684] = 3'b110;
        rom_memory[40685] = 3'b110;
        rom_memory[40686] = 3'b110;
        rom_memory[40687] = 3'b110;
        rom_memory[40688] = 3'b110;
        rom_memory[40689] = 3'b110;
        rom_memory[40690] = 3'b110;
        rom_memory[40691] = 3'b110;
        rom_memory[40692] = 3'b110;
        rom_memory[40693] = 3'b110;
        rom_memory[40694] = 3'b110;
        rom_memory[40695] = 3'b110;
        rom_memory[40696] = 3'b110;
        rom_memory[40697] = 3'b110;
        rom_memory[40698] = 3'b110;
        rom_memory[40699] = 3'b110;
        rom_memory[40700] = 3'b110;
        rom_memory[40701] = 3'b110;
        rom_memory[40702] = 3'b110;
        rom_memory[40703] = 3'b110;
        rom_memory[40704] = 3'b110;
        rom_memory[40705] = 3'b110;
        rom_memory[40706] = 3'b110;
        rom_memory[40707] = 3'b110;
        rom_memory[40708] = 3'b110;
        rom_memory[40709] = 3'b110;
        rom_memory[40710] = 3'b110;
        rom_memory[40711] = 3'b110;
        rom_memory[40712] = 3'b110;
        rom_memory[40713] = 3'b110;
        rom_memory[40714] = 3'b110;
        rom_memory[40715] = 3'b110;
        rom_memory[40716] = 3'b110;
        rom_memory[40717] = 3'b110;
        rom_memory[40718] = 3'b110;
        rom_memory[40719] = 3'b110;
        rom_memory[40720] = 3'b110;
        rom_memory[40721] = 3'b110;
        rom_memory[40722] = 3'b110;
        rom_memory[40723] = 3'b110;
        rom_memory[40724] = 3'b110;
        rom_memory[40725] = 3'b110;
        rom_memory[40726] = 3'b110;
        rom_memory[40727] = 3'b110;
        rom_memory[40728] = 3'b110;
        rom_memory[40729] = 3'b110;
        rom_memory[40730] = 3'b110;
        rom_memory[40731] = 3'b110;
        rom_memory[40732] = 3'b110;
        rom_memory[40733] = 3'b110;
        rom_memory[40734] = 3'b000;
        rom_memory[40735] = 3'b000;
        rom_memory[40736] = 3'b000;
        rom_memory[40737] = 3'b000;
        rom_memory[40738] = 3'b000;
        rom_memory[40739] = 3'b000;
        rom_memory[40740] = 3'b000;
        rom_memory[40741] = 3'b000;
        rom_memory[40742] = 3'b000;
        rom_memory[40743] = 3'b000;
        rom_memory[40744] = 3'b000;
        rom_memory[40745] = 3'b000;
        rom_memory[40746] = 3'b000;
        rom_memory[40747] = 3'b110;
        rom_memory[40748] = 3'b111;
        rom_memory[40749] = 3'b111;
        rom_memory[40750] = 3'b110;
        rom_memory[40751] = 3'b110;
        rom_memory[40752] = 3'b110;
        rom_memory[40753] = 3'b110;
        rom_memory[40754] = 3'b110;
        rom_memory[40755] = 3'b110;
        rom_memory[40756] = 3'b110;
        rom_memory[40757] = 3'b110;
        rom_memory[40758] = 3'b110;
        rom_memory[40759] = 3'b110;
        rom_memory[40760] = 3'b110;
        rom_memory[40761] = 3'b110;
        rom_memory[40762] = 3'b110;
        rom_memory[40763] = 3'b110;
        rom_memory[40764] = 3'b110;
        rom_memory[40765] = 3'b110;
        rom_memory[40766] = 3'b110;
        rom_memory[40767] = 3'b110;
        rom_memory[40768] = 3'b110;
        rom_memory[40769] = 3'b110;
        rom_memory[40770] = 3'b110;
        rom_memory[40771] = 3'b110;
        rom_memory[40772] = 3'b110;
        rom_memory[40773] = 3'b110;
        rom_memory[40774] = 3'b110;
        rom_memory[40775] = 3'b110;
        rom_memory[40776] = 3'b110;
        rom_memory[40777] = 3'b110;
        rom_memory[40778] = 3'b110;
        rom_memory[40779] = 3'b110;
        rom_memory[40780] = 3'b110;
        rom_memory[40781] = 3'b110;
        rom_memory[40782] = 3'b111;
        rom_memory[40783] = 3'b111;
        rom_memory[40784] = 3'b111;
        rom_memory[40785] = 3'b111;
        rom_memory[40786] = 3'b111;
        rom_memory[40787] = 3'b111;
        rom_memory[40788] = 3'b111;
        rom_memory[40789] = 3'b111;
        rom_memory[40790] = 3'b111;
        rom_memory[40791] = 3'b111;
        rom_memory[40792] = 3'b111;
        rom_memory[40793] = 3'b111;
        rom_memory[40794] = 3'b111;
        rom_memory[40795] = 3'b111;
        rom_memory[40796] = 3'b111;
        rom_memory[40797] = 3'b111;
        rom_memory[40798] = 3'b111;
        rom_memory[40799] = 3'b111;
        rom_memory[40800] = 3'b110;
        rom_memory[40801] = 3'b110;
        rom_memory[40802] = 3'b110;
        rom_memory[40803] = 3'b110;
        rom_memory[40804] = 3'b110;
        rom_memory[40805] = 3'b110;
        rom_memory[40806] = 3'b110;
        rom_memory[40807] = 3'b110;
        rom_memory[40808] = 3'b110;
        rom_memory[40809] = 3'b111;
        rom_memory[40810] = 3'b111;
        rom_memory[40811] = 3'b111;
        rom_memory[40812] = 3'b111;
        rom_memory[40813] = 3'b111;
        rom_memory[40814] = 3'b111;
        rom_memory[40815] = 3'b111;
        rom_memory[40816] = 3'b111;
        rom_memory[40817] = 3'b111;
        rom_memory[40818] = 3'b111;
        rom_memory[40819] = 3'b111;
        rom_memory[40820] = 3'b111;
        rom_memory[40821] = 3'b110;
        rom_memory[40822] = 3'b110;
        rom_memory[40823] = 3'b110;
        rom_memory[40824] = 3'b110;
        rom_memory[40825] = 3'b110;
        rom_memory[40826] = 3'b110;
        rom_memory[40827] = 3'b110;
        rom_memory[40828] = 3'b110;
        rom_memory[40829] = 3'b110;
        rom_memory[40830] = 3'b110;
        rom_memory[40831] = 3'b110;
        rom_memory[40832] = 3'b110;
        rom_memory[40833] = 3'b110;
        rom_memory[40834] = 3'b110;
        rom_memory[40835] = 3'b110;
        rom_memory[40836] = 3'b110;
        rom_memory[40837] = 3'b110;
        rom_memory[40838] = 3'b110;
        rom_memory[40839] = 3'b111;
        rom_memory[40840] = 3'b111;
        rom_memory[40841] = 3'b111;
        rom_memory[40842] = 3'b110;
        rom_memory[40843] = 3'b110;
        rom_memory[40844] = 3'b110;
        rom_memory[40845] = 3'b111;
        rom_memory[40846] = 3'b111;
        rom_memory[40847] = 3'b111;
        rom_memory[40848] = 3'b111;
        rom_memory[40849] = 3'b111;
        rom_memory[40850] = 3'b111;
        rom_memory[40851] = 3'b111;
        rom_memory[40852] = 3'b111;
        rom_memory[40853] = 3'b110;
        rom_memory[40854] = 3'b000;
        rom_memory[40855] = 3'b110;
        rom_memory[40856] = 3'b111;
        rom_memory[40857] = 3'b111;
        rom_memory[40858] = 3'b111;
        rom_memory[40859] = 3'b000;
        rom_memory[40860] = 3'b000;
        rom_memory[40861] = 3'b000;
        rom_memory[40862] = 3'b110;
        rom_memory[40863] = 3'b110;
        rom_memory[40864] = 3'b110;
        rom_memory[40865] = 3'b110;
        rom_memory[40866] = 3'b110;
        rom_memory[40867] = 3'b110;
        rom_memory[40868] = 3'b110;
        rom_memory[40869] = 3'b000;
        rom_memory[40870] = 3'b100;
        rom_memory[40871] = 3'b111;
        rom_memory[40872] = 3'b111;
        rom_memory[40873] = 3'b101;
        rom_memory[40874] = 3'b111;
        rom_memory[40875] = 3'b111;
        rom_memory[40876] = 3'b111;
        rom_memory[40877] = 3'b100;
        rom_memory[40878] = 3'b111;
        rom_memory[40879] = 3'b000;
        rom_memory[40880] = 3'b000;
        rom_memory[40881] = 3'b100;
        rom_memory[40882] = 3'b110;
        rom_memory[40883] = 3'b110;
        rom_memory[40884] = 3'b110;
        rom_memory[40885] = 3'b110;
        rom_memory[40886] = 3'b111;
        rom_memory[40887] = 3'b111;
        rom_memory[40888] = 3'b110;
        rom_memory[40889] = 3'b111;
        rom_memory[40890] = 3'b111;
        rom_memory[40891] = 3'b110;
        rom_memory[40892] = 3'b110;
        rom_memory[40893] = 3'b110;
        rom_memory[40894] = 3'b110;
        rom_memory[40895] = 3'b110;
        rom_memory[40896] = 3'b110;
        rom_memory[40897] = 3'b110;
        rom_memory[40898] = 3'b110;
        rom_memory[40899] = 3'b110;
        rom_memory[40900] = 3'b110;
        rom_memory[40901] = 3'b110;
        rom_memory[40902] = 3'b110;
        rom_memory[40903] = 3'b111;
        rom_memory[40904] = 3'b111;
        rom_memory[40905] = 3'b111;
        rom_memory[40906] = 3'b111;
        rom_memory[40907] = 3'b111;
        rom_memory[40908] = 3'b110;
        rom_memory[40909] = 3'b110;
        rom_memory[40910] = 3'b110;
        rom_memory[40911] = 3'b110;
        rom_memory[40912] = 3'b110;
        rom_memory[40913] = 3'b110;
        rom_memory[40914] = 3'b110;
        rom_memory[40915] = 3'b110;
        rom_memory[40916] = 3'b110;
        rom_memory[40917] = 3'b110;
        rom_memory[40918] = 3'b110;
        rom_memory[40919] = 3'b110;
        rom_memory[40920] = 3'b110;
        rom_memory[40921] = 3'b110;
        rom_memory[40922] = 3'b110;
        rom_memory[40923] = 3'b110;
        rom_memory[40924] = 3'b110;
        rom_memory[40925] = 3'b110;
        rom_memory[40926] = 3'b110;
        rom_memory[40927] = 3'b110;
        rom_memory[40928] = 3'b110;
        rom_memory[40929] = 3'b110;
        rom_memory[40930] = 3'b110;
        rom_memory[40931] = 3'b110;
        rom_memory[40932] = 3'b110;
        rom_memory[40933] = 3'b110;
        rom_memory[40934] = 3'b110;
        rom_memory[40935] = 3'b110;
        rom_memory[40936] = 3'b110;
        rom_memory[40937] = 3'b110;
        rom_memory[40938] = 3'b110;
        rom_memory[40939] = 3'b110;
        rom_memory[40940] = 3'b110;
        rom_memory[40941] = 3'b110;
        rom_memory[40942] = 3'b110;
        rom_memory[40943] = 3'b110;
        rom_memory[40944] = 3'b110;
        rom_memory[40945] = 3'b110;
        rom_memory[40946] = 3'b110;
        rom_memory[40947] = 3'b110;
        rom_memory[40948] = 3'b110;
        rom_memory[40949] = 3'b110;
        rom_memory[40950] = 3'b110;
        rom_memory[40951] = 3'b110;
        rom_memory[40952] = 3'b110;
        rom_memory[40953] = 3'b110;
        rom_memory[40954] = 3'b110;
        rom_memory[40955] = 3'b110;
        rom_memory[40956] = 3'b110;
        rom_memory[40957] = 3'b110;
        rom_memory[40958] = 3'b110;
        rom_memory[40959] = 3'b110;
        rom_memory[40960] = 3'b110;
        rom_memory[40961] = 3'b110;
        rom_memory[40962] = 3'b110;
        rom_memory[40963] = 3'b110;
        rom_memory[40964] = 3'b110;
        rom_memory[40965] = 3'b110;
        rom_memory[40966] = 3'b110;
        rom_memory[40967] = 3'b110;
        rom_memory[40968] = 3'b110;
        rom_memory[40969] = 3'b110;
        rom_memory[40970] = 3'b110;
        rom_memory[40971] = 3'b110;
        rom_memory[40972] = 3'b110;
        rom_memory[40973] = 3'b110;
        rom_memory[40974] = 3'b110;
        rom_memory[40975] = 3'b000;
        rom_memory[40976] = 3'b000;
        rom_memory[40977] = 3'b000;
        rom_memory[40978] = 3'b000;
        rom_memory[40979] = 3'b000;
        rom_memory[40980] = 3'b000;
        rom_memory[40981] = 3'b000;
        rom_memory[40982] = 3'b000;
        rom_memory[40983] = 3'b000;
        rom_memory[40984] = 3'b000;
        rom_memory[40985] = 3'b000;
        rom_memory[40986] = 3'b000;
        rom_memory[40987] = 3'b000;
        rom_memory[40988] = 3'b100;
        rom_memory[40989] = 3'b111;
        rom_memory[40990] = 3'b111;
        rom_memory[40991] = 3'b110;
        rom_memory[40992] = 3'b110;
        rom_memory[40993] = 3'b110;
        rom_memory[40994] = 3'b110;
        rom_memory[40995] = 3'b110;
        rom_memory[40996] = 3'b110;
        rom_memory[40997] = 3'b110;
        rom_memory[40998] = 3'b110;
        rom_memory[40999] = 3'b110;
        rom_memory[41000] = 3'b110;
        rom_memory[41001] = 3'b110;
        rom_memory[41002] = 3'b110;
        rom_memory[41003] = 3'b110;
        rom_memory[41004] = 3'b110;
        rom_memory[41005] = 3'b110;
        rom_memory[41006] = 3'b110;
        rom_memory[41007] = 3'b110;
        rom_memory[41008] = 3'b110;
        rom_memory[41009] = 3'b110;
        rom_memory[41010] = 3'b110;
        rom_memory[41011] = 3'b110;
        rom_memory[41012] = 3'b110;
        rom_memory[41013] = 3'b110;
        rom_memory[41014] = 3'b110;
        rom_memory[41015] = 3'b110;
        rom_memory[41016] = 3'b110;
        rom_memory[41017] = 3'b110;
        rom_memory[41018] = 3'b110;
        rom_memory[41019] = 3'b110;
        rom_memory[41020] = 3'b110;
        rom_memory[41021] = 3'b110;
        rom_memory[41022] = 3'b110;
        rom_memory[41023] = 3'b110;
        rom_memory[41024] = 3'b111;
        rom_memory[41025] = 3'b111;
        rom_memory[41026] = 3'b111;
        rom_memory[41027] = 3'b111;
        rom_memory[41028] = 3'b111;
        rom_memory[41029] = 3'b111;
        rom_memory[41030] = 3'b111;
        rom_memory[41031] = 3'b111;
        rom_memory[41032] = 3'b111;
        rom_memory[41033] = 3'b111;
        rom_memory[41034] = 3'b111;
        rom_memory[41035] = 3'b111;
        rom_memory[41036] = 3'b111;
        rom_memory[41037] = 3'b111;
        rom_memory[41038] = 3'b111;
        rom_memory[41039] = 3'b111;
        rom_memory[41040] = 3'b110;
        rom_memory[41041] = 3'b110;
        rom_memory[41042] = 3'b110;
        rom_memory[41043] = 3'b110;
        rom_memory[41044] = 3'b110;
        rom_memory[41045] = 3'b110;
        rom_memory[41046] = 3'b110;
        rom_memory[41047] = 3'b110;
        rom_memory[41048] = 3'b110;
        rom_memory[41049] = 3'b110;
        rom_memory[41050] = 3'b111;
        rom_memory[41051] = 3'b111;
        rom_memory[41052] = 3'b111;
        rom_memory[41053] = 3'b111;
        rom_memory[41054] = 3'b111;
        rom_memory[41055] = 3'b111;
        rom_memory[41056] = 3'b111;
        rom_memory[41057] = 3'b111;
        rom_memory[41058] = 3'b111;
        rom_memory[41059] = 3'b111;
        rom_memory[41060] = 3'b111;
        rom_memory[41061] = 3'b110;
        rom_memory[41062] = 3'b110;
        rom_memory[41063] = 3'b110;
        rom_memory[41064] = 3'b110;
        rom_memory[41065] = 3'b110;
        rom_memory[41066] = 3'b110;
        rom_memory[41067] = 3'b110;
        rom_memory[41068] = 3'b110;
        rom_memory[41069] = 3'b110;
        rom_memory[41070] = 3'b110;
        rom_memory[41071] = 3'b110;
        rom_memory[41072] = 3'b110;
        rom_memory[41073] = 3'b110;
        rom_memory[41074] = 3'b110;
        rom_memory[41075] = 3'b110;
        rom_memory[41076] = 3'b110;
        rom_memory[41077] = 3'b110;
        rom_memory[41078] = 3'b110;
        rom_memory[41079] = 3'b111;
        rom_memory[41080] = 3'b111;
        rom_memory[41081] = 3'b111;
        rom_memory[41082] = 3'b110;
        rom_memory[41083] = 3'b110;
        rom_memory[41084] = 3'b110;
        rom_memory[41085] = 3'b110;
        rom_memory[41086] = 3'b110;
        rom_memory[41087] = 3'b111;
        rom_memory[41088] = 3'b111;
        rom_memory[41089] = 3'b111;
        rom_memory[41090] = 3'b111;
        rom_memory[41091] = 3'b111;
        rom_memory[41092] = 3'b110;
        rom_memory[41093] = 3'b110;
        rom_memory[41094] = 3'b000;
        rom_memory[41095] = 3'b010;
        rom_memory[41096] = 3'b111;
        rom_memory[41097] = 3'b111;
        rom_memory[41098] = 3'b111;
        rom_memory[41099] = 3'b000;
        rom_memory[41100] = 3'b000;
        rom_memory[41101] = 3'b010;
        rom_memory[41102] = 3'b110;
        rom_memory[41103] = 3'b110;
        rom_memory[41104] = 3'b110;
        rom_memory[41105] = 3'b110;
        rom_memory[41106] = 3'b110;
        rom_memory[41107] = 3'b110;
        rom_memory[41108] = 3'b110;
        rom_memory[41109] = 3'b100;
        rom_memory[41110] = 3'b000;
        rom_memory[41111] = 3'b000;
        rom_memory[41112] = 3'b111;
        rom_memory[41113] = 3'b111;
        rom_memory[41114] = 3'b111;
        rom_memory[41115] = 3'b111;
        rom_memory[41116] = 3'b110;
        rom_memory[41117] = 3'b000;
        rom_memory[41118] = 3'b000;
        rom_memory[41119] = 3'b000;
        rom_memory[41120] = 3'b111;
        rom_memory[41121] = 3'b110;
        rom_memory[41122] = 3'b110;
        rom_memory[41123] = 3'b110;
        rom_memory[41124] = 3'b110;
        rom_memory[41125] = 3'b111;
        rom_memory[41126] = 3'b111;
        rom_memory[41127] = 3'b111;
        rom_memory[41128] = 3'b111;
        rom_memory[41129] = 3'b111;
        rom_memory[41130] = 3'b111;
        rom_memory[41131] = 3'b111;
        rom_memory[41132] = 3'b110;
        rom_memory[41133] = 3'b110;
        rom_memory[41134] = 3'b110;
        rom_memory[41135] = 3'b110;
        rom_memory[41136] = 3'b110;
        rom_memory[41137] = 3'b110;
        rom_memory[41138] = 3'b110;
        rom_memory[41139] = 3'b110;
        rom_memory[41140] = 3'b110;
        rom_memory[41141] = 3'b110;
        rom_memory[41142] = 3'b110;
        rom_memory[41143] = 3'b111;
        rom_memory[41144] = 3'b111;
        rom_memory[41145] = 3'b111;
        rom_memory[41146] = 3'b111;
        rom_memory[41147] = 3'b111;
        rom_memory[41148] = 3'b110;
        rom_memory[41149] = 3'b110;
        rom_memory[41150] = 3'b110;
        rom_memory[41151] = 3'b110;
        rom_memory[41152] = 3'b110;
        rom_memory[41153] = 3'b110;
        rom_memory[41154] = 3'b110;
        rom_memory[41155] = 3'b110;
        rom_memory[41156] = 3'b110;
        rom_memory[41157] = 3'b110;
        rom_memory[41158] = 3'b110;
        rom_memory[41159] = 3'b110;
        rom_memory[41160] = 3'b110;
        rom_memory[41161] = 3'b110;
        rom_memory[41162] = 3'b110;
        rom_memory[41163] = 3'b110;
        rom_memory[41164] = 3'b110;
        rom_memory[41165] = 3'b110;
        rom_memory[41166] = 3'b110;
        rom_memory[41167] = 3'b110;
        rom_memory[41168] = 3'b110;
        rom_memory[41169] = 3'b110;
        rom_memory[41170] = 3'b110;
        rom_memory[41171] = 3'b110;
        rom_memory[41172] = 3'b110;
        rom_memory[41173] = 3'b110;
        rom_memory[41174] = 3'b110;
        rom_memory[41175] = 3'b110;
        rom_memory[41176] = 3'b110;
        rom_memory[41177] = 3'b110;
        rom_memory[41178] = 3'b110;
        rom_memory[41179] = 3'b110;
        rom_memory[41180] = 3'b110;
        rom_memory[41181] = 3'b110;
        rom_memory[41182] = 3'b110;
        rom_memory[41183] = 3'b110;
        rom_memory[41184] = 3'b110;
        rom_memory[41185] = 3'b110;
        rom_memory[41186] = 3'b110;
        rom_memory[41187] = 3'b110;
        rom_memory[41188] = 3'b110;
        rom_memory[41189] = 3'b110;
        rom_memory[41190] = 3'b110;
        rom_memory[41191] = 3'b110;
        rom_memory[41192] = 3'b110;
        rom_memory[41193] = 3'b110;
        rom_memory[41194] = 3'b110;
        rom_memory[41195] = 3'b110;
        rom_memory[41196] = 3'b110;
        rom_memory[41197] = 3'b110;
        rom_memory[41198] = 3'b110;
        rom_memory[41199] = 3'b110;
        rom_memory[41200] = 3'b110;
        rom_memory[41201] = 3'b110;
        rom_memory[41202] = 3'b110;
        rom_memory[41203] = 3'b110;
        rom_memory[41204] = 3'b110;
        rom_memory[41205] = 3'b110;
        rom_memory[41206] = 3'b110;
        rom_memory[41207] = 3'b110;
        rom_memory[41208] = 3'b110;
        rom_memory[41209] = 3'b110;
        rom_memory[41210] = 3'b110;
        rom_memory[41211] = 3'b110;
        rom_memory[41212] = 3'b110;
        rom_memory[41213] = 3'b110;
        rom_memory[41214] = 3'b110;
        rom_memory[41215] = 3'b110;
        rom_memory[41216] = 3'b000;
        rom_memory[41217] = 3'b000;
        rom_memory[41218] = 3'b000;
        rom_memory[41219] = 3'b000;
        rom_memory[41220] = 3'b000;
        rom_memory[41221] = 3'b000;
        rom_memory[41222] = 3'b000;
        rom_memory[41223] = 3'b000;
        rom_memory[41224] = 3'b000;
        rom_memory[41225] = 3'b000;
        rom_memory[41226] = 3'b000;
        rom_memory[41227] = 3'b000;
        rom_memory[41228] = 3'b000;
        rom_memory[41229] = 3'b000;
        rom_memory[41230] = 3'b111;
        rom_memory[41231] = 3'b111;
        rom_memory[41232] = 3'b110;
        rom_memory[41233] = 3'b110;
        rom_memory[41234] = 3'b110;
        rom_memory[41235] = 3'b110;
        rom_memory[41236] = 3'b110;
        rom_memory[41237] = 3'b110;
        rom_memory[41238] = 3'b110;
        rom_memory[41239] = 3'b110;
        rom_memory[41240] = 3'b110;
        rom_memory[41241] = 3'b110;
        rom_memory[41242] = 3'b110;
        rom_memory[41243] = 3'b110;
        rom_memory[41244] = 3'b110;
        rom_memory[41245] = 3'b110;
        rom_memory[41246] = 3'b110;
        rom_memory[41247] = 3'b110;
        rom_memory[41248] = 3'b110;
        rom_memory[41249] = 3'b110;
        rom_memory[41250] = 3'b110;
        rom_memory[41251] = 3'b110;
        rom_memory[41252] = 3'b110;
        rom_memory[41253] = 3'b110;
        rom_memory[41254] = 3'b110;
        rom_memory[41255] = 3'b110;
        rom_memory[41256] = 3'b110;
        rom_memory[41257] = 3'b110;
        rom_memory[41258] = 3'b110;
        rom_memory[41259] = 3'b110;
        rom_memory[41260] = 3'b110;
        rom_memory[41261] = 3'b110;
        rom_memory[41262] = 3'b110;
        rom_memory[41263] = 3'b110;
        rom_memory[41264] = 3'b110;
        rom_memory[41265] = 3'b110;
        rom_memory[41266] = 3'b111;
        rom_memory[41267] = 3'b111;
        rom_memory[41268] = 3'b110;
        rom_memory[41269] = 3'b111;
        rom_memory[41270] = 3'b111;
        rom_memory[41271] = 3'b111;
        rom_memory[41272] = 3'b110;
        rom_memory[41273] = 3'b111;
        rom_memory[41274] = 3'b111;
        rom_memory[41275] = 3'b111;
        rom_memory[41276] = 3'b110;
        rom_memory[41277] = 3'b110;
        rom_memory[41278] = 3'b110;
        rom_memory[41279] = 3'b110;
        rom_memory[41280] = 3'b110;
        rom_memory[41281] = 3'b110;
        rom_memory[41282] = 3'b110;
        rom_memory[41283] = 3'b110;
        rom_memory[41284] = 3'b110;
        rom_memory[41285] = 3'b110;
        rom_memory[41286] = 3'b110;
        rom_memory[41287] = 3'b110;
        rom_memory[41288] = 3'b111;
        rom_memory[41289] = 3'b111;
        rom_memory[41290] = 3'b111;
        rom_memory[41291] = 3'b111;
        rom_memory[41292] = 3'b111;
        rom_memory[41293] = 3'b111;
        rom_memory[41294] = 3'b111;
        rom_memory[41295] = 3'b111;
        rom_memory[41296] = 3'b111;
        rom_memory[41297] = 3'b111;
        rom_memory[41298] = 3'b111;
        rom_memory[41299] = 3'b110;
        rom_memory[41300] = 3'b110;
        rom_memory[41301] = 3'b110;
        rom_memory[41302] = 3'b110;
        rom_memory[41303] = 3'b110;
        rom_memory[41304] = 3'b110;
        rom_memory[41305] = 3'b110;
        rom_memory[41306] = 3'b110;
        rom_memory[41307] = 3'b110;
        rom_memory[41308] = 3'b110;
        rom_memory[41309] = 3'b110;
        rom_memory[41310] = 3'b110;
        rom_memory[41311] = 3'b110;
        rom_memory[41312] = 3'b110;
        rom_memory[41313] = 3'b110;
        rom_memory[41314] = 3'b110;
        rom_memory[41315] = 3'b110;
        rom_memory[41316] = 3'b110;
        rom_memory[41317] = 3'b110;
        rom_memory[41318] = 3'b111;
        rom_memory[41319] = 3'b111;
        rom_memory[41320] = 3'b111;
        rom_memory[41321] = 3'b111;
        rom_memory[41322] = 3'b111;
        rom_memory[41323] = 3'b110;
        rom_memory[41324] = 3'b110;
        rom_memory[41325] = 3'b110;
        rom_memory[41326] = 3'b110;
        rom_memory[41327] = 3'b110;
        rom_memory[41328] = 3'b110;
        rom_memory[41329] = 3'b111;
        rom_memory[41330] = 3'b111;
        rom_memory[41331] = 3'b111;
        rom_memory[41332] = 3'b110;
        rom_memory[41333] = 3'b110;
        rom_memory[41334] = 3'b000;
        rom_memory[41335] = 3'b111;
        rom_memory[41336] = 3'b111;
        rom_memory[41337] = 3'b111;
        rom_memory[41338] = 3'b111;
        rom_memory[41339] = 3'b000;
        rom_memory[41340] = 3'b010;
        rom_memory[41341] = 3'b111;
        rom_memory[41342] = 3'b110;
        rom_memory[41343] = 3'b110;
        rom_memory[41344] = 3'b110;
        rom_memory[41345] = 3'b110;
        rom_memory[41346] = 3'b110;
        rom_memory[41347] = 3'b110;
        rom_memory[41348] = 3'b110;
        rom_memory[41349] = 3'b110;
        rom_memory[41350] = 3'b110;
        rom_memory[41351] = 3'b100;
        rom_memory[41352] = 3'b100;
        rom_memory[41353] = 3'b111;
        rom_memory[41354] = 3'b111;
        rom_memory[41355] = 3'b110;
        rom_memory[41356] = 3'b110;
        rom_memory[41357] = 3'b000;
        rom_memory[41358] = 3'b000;
        rom_memory[41359] = 3'b100;
        rom_memory[41360] = 3'b111;
        rom_memory[41361] = 3'b110;
        rom_memory[41362] = 3'b110;
        rom_memory[41363] = 3'b110;
        rom_memory[41364] = 3'b111;
        rom_memory[41365] = 3'b111;
        rom_memory[41366] = 3'b111;
        rom_memory[41367] = 3'b111;
        rom_memory[41368] = 3'b111;
        rom_memory[41369] = 3'b111;
        rom_memory[41370] = 3'b111;
        rom_memory[41371] = 3'b110;
        rom_memory[41372] = 3'b110;
        rom_memory[41373] = 3'b110;
        rom_memory[41374] = 3'b110;
        rom_memory[41375] = 3'b110;
        rom_memory[41376] = 3'b110;
        rom_memory[41377] = 3'b110;
        rom_memory[41378] = 3'b110;
        rom_memory[41379] = 3'b110;
        rom_memory[41380] = 3'b110;
        rom_memory[41381] = 3'b110;
        rom_memory[41382] = 3'b110;
        rom_memory[41383] = 3'b111;
        rom_memory[41384] = 3'b111;
        rom_memory[41385] = 3'b111;
        rom_memory[41386] = 3'b111;
        rom_memory[41387] = 3'b111;
        rom_memory[41388] = 3'b110;
        rom_memory[41389] = 3'b110;
        rom_memory[41390] = 3'b110;
        rom_memory[41391] = 3'b110;
        rom_memory[41392] = 3'b110;
        rom_memory[41393] = 3'b110;
        rom_memory[41394] = 3'b110;
        rom_memory[41395] = 3'b110;
        rom_memory[41396] = 3'b110;
        rom_memory[41397] = 3'b110;
        rom_memory[41398] = 3'b110;
        rom_memory[41399] = 3'b110;
        rom_memory[41400] = 3'b110;
        rom_memory[41401] = 3'b110;
        rom_memory[41402] = 3'b110;
        rom_memory[41403] = 3'b110;
        rom_memory[41404] = 3'b110;
        rom_memory[41405] = 3'b110;
        rom_memory[41406] = 3'b110;
        rom_memory[41407] = 3'b110;
        rom_memory[41408] = 3'b110;
        rom_memory[41409] = 3'b110;
        rom_memory[41410] = 3'b110;
        rom_memory[41411] = 3'b110;
        rom_memory[41412] = 3'b110;
        rom_memory[41413] = 3'b110;
        rom_memory[41414] = 3'b110;
        rom_memory[41415] = 3'b110;
        rom_memory[41416] = 3'b110;
        rom_memory[41417] = 3'b110;
        rom_memory[41418] = 3'b110;
        rom_memory[41419] = 3'b110;
        rom_memory[41420] = 3'b110;
        rom_memory[41421] = 3'b110;
        rom_memory[41422] = 3'b110;
        rom_memory[41423] = 3'b110;
        rom_memory[41424] = 3'b110;
        rom_memory[41425] = 3'b110;
        rom_memory[41426] = 3'b110;
        rom_memory[41427] = 3'b110;
        rom_memory[41428] = 3'b110;
        rom_memory[41429] = 3'b110;
        rom_memory[41430] = 3'b110;
        rom_memory[41431] = 3'b110;
        rom_memory[41432] = 3'b110;
        rom_memory[41433] = 3'b110;
        rom_memory[41434] = 3'b110;
        rom_memory[41435] = 3'b110;
        rom_memory[41436] = 3'b110;
        rom_memory[41437] = 3'b110;
        rom_memory[41438] = 3'b110;
        rom_memory[41439] = 3'b110;
        rom_memory[41440] = 3'b110;
        rom_memory[41441] = 3'b110;
        rom_memory[41442] = 3'b110;
        rom_memory[41443] = 3'b110;
        rom_memory[41444] = 3'b110;
        rom_memory[41445] = 3'b110;
        rom_memory[41446] = 3'b110;
        rom_memory[41447] = 3'b110;
        rom_memory[41448] = 3'b110;
        rom_memory[41449] = 3'b110;
        rom_memory[41450] = 3'b110;
        rom_memory[41451] = 3'b110;
        rom_memory[41452] = 3'b110;
        rom_memory[41453] = 3'b110;
        rom_memory[41454] = 3'b110;
        rom_memory[41455] = 3'b110;
        rom_memory[41456] = 3'b110;
        rom_memory[41457] = 3'b000;
        rom_memory[41458] = 3'b000;
        rom_memory[41459] = 3'b000;
        rom_memory[41460] = 3'b000;
        rom_memory[41461] = 3'b000;
        rom_memory[41462] = 3'b000;
        rom_memory[41463] = 3'b000;
        rom_memory[41464] = 3'b000;
        rom_memory[41465] = 3'b000;
        rom_memory[41466] = 3'b000;
        rom_memory[41467] = 3'b000;
        rom_memory[41468] = 3'b000;
        rom_memory[41469] = 3'b000;
        rom_memory[41470] = 3'b000;
        rom_memory[41471] = 3'b110;
        rom_memory[41472] = 3'b111;
        rom_memory[41473] = 3'b111;
        rom_memory[41474] = 3'b110;
        rom_memory[41475] = 3'b110;
        rom_memory[41476] = 3'b110;
        rom_memory[41477] = 3'b110;
        rom_memory[41478] = 3'b110;
        rom_memory[41479] = 3'b110;
        rom_memory[41480] = 3'b110;
        rom_memory[41481] = 3'b110;
        rom_memory[41482] = 3'b110;
        rom_memory[41483] = 3'b110;
        rom_memory[41484] = 3'b110;
        rom_memory[41485] = 3'b110;
        rom_memory[41486] = 3'b110;
        rom_memory[41487] = 3'b110;
        rom_memory[41488] = 3'b110;
        rom_memory[41489] = 3'b110;
        rom_memory[41490] = 3'b110;
        rom_memory[41491] = 3'b110;
        rom_memory[41492] = 3'b110;
        rom_memory[41493] = 3'b110;
        rom_memory[41494] = 3'b110;
        rom_memory[41495] = 3'b110;
        rom_memory[41496] = 3'b110;
        rom_memory[41497] = 3'b110;
        rom_memory[41498] = 3'b110;
        rom_memory[41499] = 3'b110;
        rom_memory[41500] = 3'b110;
        rom_memory[41501] = 3'b110;
        rom_memory[41502] = 3'b110;
        rom_memory[41503] = 3'b110;
        rom_memory[41504] = 3'b110;
        rom_memory[41505] = 3'b110;
        rom_memory[41506] = 3'b110;
        rom_memory[41507] = 3'b111;
        rom_memory[41508] = 3'b110;
        rom_memory[41509] = 3'b111;
        rom_memory[41510] = 3'b111;
        rom_memory[41511] = 3'b110;
        rom_memory[41512] = 3'b110;
        rom_memory[41513] = 3'b111;
        rom_memory[41514] = 3'b111;
        rom_memory[41515] = 3'b111;
        rom_memory[41516] = 3'b110;
        rom_memory[41517] = 3'b110;
        rom_memory[41518] = 3'b110;
        rom_memory[41519] = 3'b110;
        rom_memory[41520] = 3'b110;
        rom_memory[41521] = 3'b110;
        rom_memory[41522] = 3'b110;
        rom_memory[41523] = 3'b110;
        rom_memory[41524] = 3'b110;
        rom_memory[41525] = 3'b110;
        rom_memory[41526] = 3'b110;
        rom_memory[41527] = 3'b111;
        rom_memory[41528] = 3'b111;
        rom_memory[41529] = 3'b111;
        rom_memory[41530] = 3'b111;
        rom_memory[41531] = 3'b111;
        rom_memory[41532] = 3'b111;
        rom_memory[41533] = 3'b111;
        rom_memory[41534] = 3'b111;
        rom_memory[41535] = 3'b111;
        rom_memory[41536] = 3'b111;
        rom_memory[41537] = 3'b111;
        rom_memory[41538] = 3'b111;
        rom_memory[41539] = 3'b111;
        rom_memory[41540] = 3'b110;
        rom_memory[41541] = 3'b110;
        rom_memory[41542] = 3'b110;
        rom_memory[41543] = 3'b110;
        rom_memory[41544] = 3'b110;
        rom_memory[41545] = 3'b110;
        rom_memory[41546] = 3'b110;
        rom_memory[41547] = 3'b110;
        rom_memory[41548] = 3'b110;
        rom_memory[41549] = 3'b110;
        rom_memory[41550] = 3'b110;
        rom_memory[41551] = 3'b110;
        rom_memory[41552] = 3'b110;
        rom_memory[41553] = 3'b110;
        rom_memory[41554] = 3'b110;
        rom_memory[41555] = 3'b110;
        rom_memory[41556] = 3'b111;
        rom_memory[41557] = 3'b111;
        rom_memory[41558] = 3'b111;
        rom_memory[41559] = 3'b111;
        rom_memory[41560] = 3'b111;
        rom_memory[41561] = 3'b111;
        rom_memory[41562] = 3'b111;
        rom_memory[41563] = 3'b111;
        rom_memory[41564] = 3'b110;
        rom_memory[41565] = 3'b110;
        rom_memory[41566] = 3'b110;
        rom_memory[41567] = 3'b110;
        rom_memory[41568] = 3'b110;
        rom_memory[41569] = 3'b110;
        rom_memory[41570] = 3'b110;
        rom_memory[41571] = 3'b111;
        rom_memory[41572] = 3'b111;
        rom_memory[41573] = 3'b110;
        rom_memory[41574] = 3'b110;
        rom_memory[41575] = 3'b111;
        rom_memory[41576] = 3'b111;
        rom_memory[41577] = 3'b111;
        rom_memory[41578] = 3'b110;
        rom_memory[41579] = 3'b000;
        rom_memory[41580] = 3'b110;
        rom_memory[41581] = 3'b111;
        rom_memory[41582] = 3'b110;
        rom_memory[41583] = 3'b110;
        rom_memory[41584] = 3'b110;
        rom_memory[41585] = 3'b110;
        rom_memory[41586] = 3'b110;
        rom_memory[41587] = 3'b110;
        rom_memory[41588] = 3'b110;
        rom_memory[41589] = 3'b110;
        rom_memory[41590] = 3'b111;
        rom_memory[41591] = 3'b110;
        rom_memory[41592] = 3'b100;
        rom_memory[41593] = 3'b111;
        rom_memory[41594] = 3'b111;
        rom_memory[41595] = 3'b111;
        rom_memory[41596] = 3'b000;
        rom_memory[41597] = 3'b000;
        rom_memory[41598] = 3'b111;
        rom_memory[41599] = 3'b100;
        rom_memory[41600] = 3'b110;
        rom_memory[41601] = 3'b110;
        rom_memory[41602] = 3'b110;
        rom_memory[41603] = 3'b111;
        rom_memory[41604] = 3'b111;
        rom_memory[41605] = 3'b111;
        rom_memory[41606] = 3'b111;
        rom_memory[41607] = 3'b111;
        rom_memory[41608] = 3'b111;
        rom_memory[41609] = 3'b111;
        rom_memory[41610] = 3'b111;
        rom_memory[41611] = 3'b111;
        rom_memory[41612] = 3'b111;
        rom_memory[41613] = 3'b110;
        rom_memory[41614] = 3'b110;
        rom_memory[41615] = 3'b110;
        rom_memory[41616] = 3'b110;
        rom_memory[41617] = 3'b110;
        rom_memory[41618] = 3'b110;
        rom_memory[41619] = 3'b110;
        rom_memory[41620] = 3'b110;
        rom_memory[41621] = 3'b110;
        rom_memory[41622] = 3'b110;
        rom_memory[41623] = 3'b111;
        rom_memory[41624] = 3'b111;
        rom_memory[41625] = 3'b111;
        rom_memory[41626] = 3'b111;
        rom_memory[41627] = 3'b111;
        rom_memory[41628] = 3'b111;
        rom_memory[41629] = 3'b110;
        rom_memory[41630] = 3'b110;
        rom_memory[41631] = 3'b110;
        rom_memory[41632] = 3'b110;
        rom_memory[41633] = 3'b110;
        rom_memory[41634] = 3'b110;
        rom_memory[41635] = 3'b110;
        rom_memory[41636] = 3'b110;
        rom_memory[41637] = 3'b110;
        rom_memory[41638] = 3'b110;
        rom_memory[41639] = 3'b110;
        rom_memory[41640] = 3'b110;
        rom_memory[41641] = 3'b110;
        rom_memory[41642] = 3'b110;
        rom_memory[41643] = 3'b110;
        rom_memory[41644] = 3'b110;
        rom_memory[41645] = 3'b110;
        rom_memory[41646] = 3'b110;
        rom_memory[41647] = 3'b110;
        rom_memory[41648] = 3'b110;
        rom_memory[41649] = 3'b110;
        rom_memory[41650] = 3'b110;
        rom_memory[41651] = 3'b110;
        rom_memory[41652] = 3'b110;
        rom_memory[41653] = 3'b110;
        rom_memory[41654] = 3'b110;
        rom_memory[41655] = 3'b110;
        rom_memory[41656] = 3'b110;
        rom_memory[41657] = 3'b110;
        rom_memory[41658] = 3'b110;
        rom_memory[41659] = 3'b110;
        rom_memory[41660] = 3'b110;
        rom_memory[41661] = 3'b110;
        rom_memory[41662] = 3'b110;
        rom_memory[41663] = 3'b110;
        rom_memory[41664] = 3'b110;
        rom_memory[41665] = 3'b110;
        rom_memory[41666] = 3'b110;
        rom_memory[41667] = 3'b110;
        rom_memory[41668] = 3'b110;
        rom_memory[41669] = 3'b110;
        rom_memory[41670] = 3'b110;
        rom_memory[41671] = 3'b110;
        rom_memory[41672] = 3'b110;
        rom_memory[41673] = 3'b110;
        rom_memory[41674] = 3'b110;
        rom_memory[41675] = 3'b110;
        rom_memory[41676] = 3'b110;
        rom_memory[41677] = 3'b110;
        rom_memory[41678] = 3'b110;
        rom_memory[41679] = 3'b110;
        rom_memory[41680] = 3'b110;
        rom_memory[41681] = 3'b110;
        rom_memory[41682] = 3'b110;
        rom_memory[41683] = 3'b110;
        rom_memory[41684] = 3'b110;
        rom_memory[41685] = 3'b110;
        rom_memory[41686] = 3'b110;
        rom_memory[41687] = 3'b110;
        rom_memory[41688] = 3'b110;
        rom_memory[41689] = 3'b110;
        rom_memory[41690] = 3'b110;
        rom_memory[41691] = 3'b110;
        rom_memory[41692] = 3'b110;
        rom_memory[41693] = 3'b110;
        rom_memory[41694] = 3'b110;
        rom_memory[41695] = 3'b110;
        rom_memory[41696] = 3'b110;
        rom_memory[41697] = 3'b110;
        rom_memory[41698] = 3'b100;
        rom_memory[41699] = 3'b000;
        rom_memory[41700] = 3'b000;
        rom_memory[41701] = 3'b000;
        rom_memory[41702] = 3'b000;
        rom_memory[41703] = 3'b000;
        rom_memory[41704] = 3'b000;
        rom_memory[41705] = 3'b000;
        rom_memory[41706] = 3'b000;
        rom_memory[41707] = 3'b000;
        rom_memory[41708] = 3'b000;
        rom_memory[41709] = 3'b000;
        rom_memory[41710] = 3'b000;
        rom_memory[41711] = 3'b000;
        rom_memory[41712] = 3'b000;
        rom_memory[41713] = 3'b111;
        rom_memory[41714] = 3'b111;
        rom_memory[41715] = 3'b110;
        rom_memory[41716] = 3'b110;
        rom_memory[41717] = 3'b110;
        rom_memory[41718] = 3'b110;
        rom_memory[41719] = 3'b110;
        rom_memory[41720] = 3'b110;
        rom_memory[41721] = 3'b110;
        rom_memory[41722] = 3'b110;
        rom_memory[41723] = 3'b110;
        rom_memory[41724] = 3'b110;
        rom_memory[41725] = 3'b110;
        rom_memory[41726] = 3'b110;
        rom_memory[41727] = 3'b110;
        rom_memory[41728] = 3'b110;
        rom_memory[41729] = 3'b110;
        rom_memory[41730] = 3'b110;
        rom_memory[41731] = 3'b110;
        rom_memory[41732] = 3'b110;
        rom_memory[41733] = 3'b110;
        rom_memory[41734] = 3'b110;
        rom_memory[41735] = 3'b110;
        rom_memory[41736] = 3'b110;
        rom_memory[41737] = 3'b110;
        rom_memory[41738] = 3'b110;
        rom_memory[41739] = 3'b110;
        rom_memory[41740] = 3'b110;
        rom_memory[41741] = 3'b110;
        rom_memory[41742] = 3'b110;
        rom_memory[41743] = 3'b110;
        rom_memory[41744] = 3'b110;
        rom_memory[41745] = 3'b110;
        rom_memory[41746] = 3'b110;
        rom_memory[41747] = 3'b110;
        rom_memory[41748] = 3'b110;
        rom_memory[41749] = 3'b110;
        rom_memory[41750] = 3'b110;
        rom_memory[41751] = 3'b110;
        rom_memory[41752] = 3'b110;
        rom_memory[41753] = 3'b110;
        rom_memory[41754] = 3'b110;
        rom_memory[41755] = 3'b110;
        rom_memory[41756] = 3'b110;
        rom_memory[41757] = 3'b110;
        rom_memory[41758] = 3'b110;
        rom_memory[41759] = 3'b110;
        rom_memory[41760] = 3'b110;
        rom_memory[41761] = 3'b110;
        rom_memory[41762] = 3'b110;
        rom_memory[41763] = 3'b110;
        rom_memory[41764] = 3'b110;
        rom_memory[41765] = 3'b110;
        rom_memory[41766] = 3'b110;
        rom_memory[41767] = 3'b111;
        rom_memory[41768] = 3'b111;
        rom_memory[41769] = 3'b111;
        rom_memory[41770] = 3'b111;
        rom_memory[41771] = 3'b111;
        rom_memory[41772] = 3'b111;
        rom_memory[41773] = 3'b111;
        rom_memory[41774] = 3'b111;
        rom_memory[41775] = 3'b111;
        rom_memory[41776] = 3'b111;
        rom_memory[41777] = 3'b111;
        rom_memory[41778] = 3'b111;
        rom_memory[41779] = 3'b110;
        rom_memory[41780] = 3'b110;
        rom_memory[41781] = 3'b110;
        rom_memory[41782] = 3'b110;
        rom_memory[41783] = 3'b110;
        rom_memory[41784] = 3'b110;
        rom_memory[41785] = 3'b110;
        rom_memory[41786] = 3'b110;
        rom_memory[41787] = 3'b110;
        rom_memory[41788] = 3'b110;
        rom_memory[41789] = 3'b110;
        rom_memory[41790] = 3'b110;
        rom_memory[41791] = 3'b110;
        rom_memory[41792] = 3'b110;
        rom_memory[41793] = 3'b110;
        rom_memory[41794] = 3'b110;
        rom_memory[41795] = 3'b110;
        rom_memory[41796] = 3'b111;
        rom_memory[41797] = 3'b111;
        rom_memory[41798] = 3'b111;
        rom_memory[41799] = 3'b111;
        rom_memory[41800] = 3'b111;
        rom_memory[41801] = 3'b111;
        rom_memory[41802] = 3'b111;
        rom_memory[41803] = 3'b111;
        rom_memory[41804] = 3'b111;
        rom_memory[41805] = 3'b110;
        rom_memory[41806] = 3'b110;
        rom_memory[41807] = 3'b110;
        rom_memory[41808] = 3'b110;
        rom_memory[41809] = 3'b110;
        rom_memory[41810] = 3'b110;
        rom_memory[41811] = 3'b110;
        rom_memory[41812] = 3'b111;
        rom_memory[41813] = 3'b110;
        rom_memory[41814] = 3'b110;
        rom_memory[41815] = 3'b111;
        rom_memory[41816] = 3'b111;
        rom_memory[41817] = 3'b111;
        rom_memory[41818] = 3'b110;
        rom_memory[41819] = 3'b100;
        rom_memory[41820] = 3'b110;
        rom_memory[41821] = 3'b111;
        rom_memory[41822] = 3'b111;
        rom_memory[41823] = 3'b110;
        rom_memory[41824] = 3'b110;
        rom_memory[41825] = 3'b110;
        rom_memory[41826] = 3'b110;
        rom_memory[41827] = 3'b110;
        rom_memory[41828] = 3'b110;
        rom_memory[41829] = 3'b110;
        rom_memory[41830] = 3'b111;
        rom_memory[41831] = 3'b111;
        rom_memory[41832] = 3'b100;
        rom_memory[41833] = 3'b100;
        rom_memory[41834] = 3'b111;
        rom_memory[41835] = 3'b111;
        rom_memory[41836] = 3'b000;
        rom_memory[41837] = 3'b000;
        rom_memory[41838] = 3'b000;
        rom_memory[41839] = 3'b100;
        rom_memory[41840] = 3'b110;
        rom_memory[41841] = 3'b111;
        rom_memory[41842] = 3'b111;
        rom_memory[41843] = 3'b111;
        rom_memory[41844] = 3'b111;
        rom_memory[41845] = 3'b111;
        rom_memory[41846] = 3'b111;
        rom_memory[41847] = 3'b111;
        rom_memory[41848] = 3'b111;
        rom_memory[41849] = 3'b111;
        rom_memory[41850] = 3'b111;
        rom_memory[41851] = 3'b111;
        rom_memory[41852] = 3'b111;
        rom_memory[41853] = 3'b111;
        rom_memory[41854] = 3'b110;
        rom_memory[41855] = 3'b110;
        rom_memory[41856] = 3'b110;
        rom_memory[41857] = 3'b110;
        rom_memory[41858] = 3'b110;
        rom_memory[41859] = 3'b110;
        rom_memory[41860] = 3'b110;
        rom_memory[41861] = 3'b110;
        rom_memory[41862] = 3'b110;
        rom_memory[41863] = 3'b111;
        rom_memory[41864] = 3'b111;
        rom_memory[41865] = 3'b111;
        rom_memory[41866] = 3'b111;
        rom_memory[41867] = 3'b111;
        rom_memory[41868] = 3'b111;
        rom_memory[41869] = 3'b111;
        rom_memory[41870] = 3'b110;
        rom_memory[41871] = 3'b110;
        rom_memory[41872] = 3'b110;
        rom_memory[41873] = 3'b110;
        rom_memory[41874] = 3'b110;
        rom_memory[41875] = 3'b110;
        rom_memory[41876] = 3'b110;
        rom_memory[41877] = 3'b110;
        rom_memory[41878] = 3'b110;
        rom_memory[41879] = 3'b110;
        rom_memory[41880] = 3'b110;
        rom_memory[41881] = 3'b110;
        rom_memory[41882] = 3'b110;
        rom_memory[41883] = 3'b110;
        rom_memory[41884] = 3'b110;
        rom_memory[41885] = 3'b110;
        rom_memory[41886] = 3'b110;
        rom_memory[41887] = 3'b110;
        rom_memory[41888] = 3'b110;
        rom_memory[41889] = 3'b110;
        rom_memory[41890] = 3'b110;
        rom_memory[41891] = 3'b110;
        rom_memory[41892] = 3'b110;
        rom_memory[41893] = 3'b110;
        rom_memory[41894] = 3'b110;
        rom_memory[41895] = 3'b110;
        rom_memory[41896] = 3'b110;
        rom_memory[41897] = 3'b110;
        rom_memory[41898] = 3'b110;
        rom_memory[41899] = 3'b110;
        rom_memory[41900] = 3'b110;
        rom_memory[41901] = 3'b110;
        rom_memory[41902] = 3'b110;
        rom_memory[41903] = 3'b110;
        rom_memory[41904] = 3'b110;
        rom_memory[41905] = 3'b110;
        rom_memory[41906] = 3'b110;
        rom_memory[41907] = 3'b110;
        rom_memory[41908] = 3'b110;
        rom_memory[41909] = 3'b110;
        rom_memory[41910] = 3'b110;
        rom_memory[41911] = 3'b110;
        rom_memory[41912] = 3'b110;
        rom_memory[41913] = 3'b110;
        rom_memory[41914] = 3'b110;
        rom_memory[41915] = 3'b110;
        rom_memory[41916] = 3'b110;
        rom_memory[41917] = 3'b110;
        rom_memory[41918] = 3'b110;
        rom_memory[41919] = 3'b110;
        rom_memory[41920] = 3'b110;
        rom_memory[41921] = 3'b110;
        rom_memory[41922] = 3'b110;
        rom_memory[41923] = 3'b110;
        rom_memory[41924] = 3'b110;
        rom_memory[41925] = 3'b110;
        rom_memory[41926] = 3'b110;
        rom_memory[41927] = 3'b110;
        rom_memory[41928] = 3'b110;
        rom_memory[41929] = 3'b110;
        rom_memory[41930] = 3'b110;
        rom_memory[41931] = 3'b110;
        rom_memory[41932] = 3'b110;
        rom_memory[41933] = 3'b110;
        rom_memory[41934] = 3'b110;
        rom_memory[41935] = 3'b110;
        rom_memory[41936] = 3'b110;
        rom_memory[41937] = 3'b110;
        rom_memory[41938] = 3'b110;
        rom_memory[41939] = 3'b110;
        rom_memory[41940] = 3'b000;
        rom_memory[41941] = 3'b000;
        rom_memory[41942] = 3'b000;
        rom_memory[41943] = 3'b000;
        rom_memory[41944] = 3'b000;
        rom_memory[41945] = 3'b000;
        rom_memory[41946] = 3'b000;
        rom_memory[41947] = 3'b000;
        rom_memory[41948] = 3'b000;
        rom_memory[41949] = 3'b000;
        rom_memory[41950] = 3'b000;
        rom_memory[41951] = 3'b000;
        rom_memory[41952] = 3'b000;
        rom_memory[41953] = 3'b000;
        rom_memory[41954] = 3'b110;
        rom_memory[41955] = 3'b111;
        rom_memory[41956] = 3'b110;
        rom_memory[41957] = 3'b110;
        rom_memory[41958] = 3'b110;
        rom_memory[41959] = 3'b110;
        rom_memory[41960] = 3'b110;
        rom_memory[41961] = 3'b110;
        rom_memory[41962] = 3'b110;
        rom_memory[41963] = 3'b110;
        rom_memory[41964] = 3'b110;
        rom_memory[41965] = 3'b110;
        rom_memory[41966] = 3'b110;
        rom_memory[41967] = 3'b110;
        rom_memory[41968] = 3'b110;
        rom_memory[41969] = 3'b110;
        rom_memory[41970] = 3'b110;
        rom_memory[41971] = 3'b110;
        rom_memory[41972] = 3'b110;
        rom_memory[41973] = 3'b110;
        rom_memory[41974] = 3'b110;
        rom_memory[41975] = 3'b110;
        rom_memory[41976] = 3'b110;
        rom_memory[41977] = 3'b110;
        rom_memory[41978] = 3'b110;
        rom_memory[41979] = 3'b110;
        rom_memory[41980] = 3'b110;
        rom_memory[41981] = 3'b110;
        rom_memory[41982] = 3'b110;
        rom_memory[41983] = 3'b110;
        rom_memory[41984] = 3'b110;
        rom_memory[41985] = 3'b110;
        rom_memory[41986] = 3'b110;
        rom_memory[41987] = 3'b110;
        rom_memory[41988] = 3'b110;
        rom_memory[41989] = 3'b110;
        rom_memory[41990] = 3'b110;
        rom_memory[41991] = 3'b110;
        rom_memory[41992] = 3'b110;
        rom_memory[41993] = 3'b110;
        rom_memory[41994] = 3'b110;
        rom_memory[41995] = 3'b110;
        rom_memory[41996] = 3'b110;
        rom_memory[41997] = 3'b110;
        rom_memory[41998] = 3'b110;
        rom_memory[41999] = 3'b110;
        rom_memory[42000] = 3'b110;
        rom_memory[42001] = 3'b110;
        rom_memory[42002] = 3'b110;
        rom_memory[42003] = 3'b110;
        rom_memory[42004] = 3'b110;
        rom_memory[42005] = 3'b110;
        rom_memory[42006] = 3'b111;
        rom_memory[42007] = 3'b111;
        rom_memory[42008] = 3'b111;
        rom_memory[42009] = 3'b111;
        rom_memory[42010] = 3'b111;
        rom_memory[42011] = 3'b111;
        rom_memory[42012] = 3'b111;
        rom_memory[42013] = 3'b111;
        rom_memory[42014] = 3'b111;
        rom_memory[42015] = 3'b111;
        rom_memory[42016] = 3'b111;
        rom_memory[42017] = 3'b111;
        rom_memory[42018] = 3'b111;
        rom_memory[42019] = 3'b111;
        rom_memory[42020] = 3'b110;
        rom_memory[42021] = 3'b110;
        rom_memory[42022] = 3'b110;
        rom_memory[42023] = 3'b110;
        rom_memory[42024] = 3'b110;
        rom_memory[42025] = 3'b110;
        rom_memory[42026] = 3'b110;
        rom_memory[42027] = 3'b110;
        rom_memory[42028] = 3'b110;
        rom_memory[42029] = 3'b110;
        rom_memory[42030] = 3'b110;
        rom_memory[42031] = 3'b110;
        rom_memory[42032] = 3'b110;
        rom_memory[42033] = 3'b110;
        rom_memory[42034] = 3'b110;
        rom_memory[42035] = 3'b110;
        rom_memory[42036] = 3'b110;
        rom_memory[42037] = 3'b111;
        rom_memory[42038] = 3'b111;
        rom_memory[42039] = 3'b111;
        rom_memory[42040] = 3'b111;
        rom_memory[42041] = 3'b111;
        rom_memory[42042] = 3'b111;
        rom_memory[42043] = 3'b110;
        rom_memory[42044] = 3'b111;
        rom_memory[42045] = 3'b111;
        rom_memory[42046] = 3'b110;
        rom_memory[42047] = 3'b110;
        rom_memory[42048] = 3'b110;
        rom_memory[42049] = 3'b110;
        rom_memory[42050] = 3'b110;
        rom_memory[42051] = 3'b110;
        rom_memory[42052] = 3'b111;
        rom_memory[42053] = 3'b111;
        rom_memory[42054] = 3'b111;
        rom_memory[42055] = 3'b111;
        rom_memory[42056] = 3'b111;
        rom_memory[42057] = 3'b111;
        rom_memory[42058] = 3'b110;
        rom_memory[42059] = 3'b100;
        rom_memory[42060] = 3'b110;
        rom_memory[42061] = 3'b110;
        rom_memory[42062] = 3'b111;
        rom_memory[42063] = 3'b110;
        rom_memory[42064] = 3'b110;
        rom_memory[42065] = 3'b110;
        rom_memory[42066] = 3'b110;
        rom_memory[42067] = 3'b110;
        rom_memory[42068] = 3'b110;
        rom_memory[42069] = 3'b111;
        rom_memory[42070] = 3'b111;
        rom_memory[42071] = 3'b111;
        rom_memory[42072] = 3'b100;
        rom_memory[42073] = 3'b100;
        rom_memory[42074] = 3'b100;
        rom_memory[42075] = 3'b111;
        rom_memory[42076] = 3'b000;
        rom_memory[42077] = 3'b110;
        rom_memory[42078] = 3'b111;
        rom_memory[42079] = 3'b111;
        rom_memory[42080] = 3'b110;
        rom_memory[42081] = 3'b111;
        rom_memory[42082] = 3'b111;
        rom_memory[42083] = 3'b111;
        rom_memory[42084] = 3'b111;
        rom_memory[42085] = 3'b111;
        rom_memory[42086] = 3'b111;
        rom_memory[42087] = 3'b111;
        rom_memory[42088] = 3'b111;
        rom_memory[42089] = 3'b111;
        rom_memory[42090] = 3'b111;
        rom_memory[42091] = 3'b111;
        rom_memory[42092] = 3'b111;
        rom_memory[42093] = 3'b111;
        rom_memory[42094] = 3'b110;
        rom_memory[42095] = 3'b110;
        rom_memory[42096] = 3'b110;
        rom_memory[42097] = 3'b110;
        rom_memory[42098] = 3'b110;
        rom_memory[42099] = 3'b110;
        rom_memory[42100] = 3'b110;
        rom_memory[42101] = 3'b110;
        rom_memory[42102] = 3'b111;
        rom_memory[42103] = 3'b111;
        rom_memory[42104] = 3'b111;
        rom_memory[42105] = 3'b111;
        rom_memory[42106] = 3'b111;
        rom_memory[42107] = 3'b111;
        rom_memory[42108] = 3'b111;
        rom_memory[42109] = 3'b111;
        rom_memory[42110] = 3'b111;
        rom_memory[42111] = 3'b110;
        rom_memory[42112] = 3'b110;
        rom_memory[42113] = 3'b110;
        rom_memory[42114] = 3'b110;
        rom_memory[42115] = 3'b110;
        rom_memory[42116] = 3'b110;
        rom_memory[42117] = 3'b110;
        rom_memory[42118] = 3'b110;
        rom_memory[42119] = 3'b110;
        rom_memory[42120] = 3'b110;
        rom_memory[42121] = 3'b110;
        rom_memory[42122] = 3'b110;
        rom_memory[42123] = 3'b110;
        rom_memory[42124] = 3'b110;
        rom_memory[42125] = 3'b110;
        rom_memory[42126] = 3'b110;
        rom_memory[42127] = 3'b110;
        rom_memory[42128] = 3'b110;
        rom_memory[42129] = 3'b110;
        rom_memory[42130] = 3'b110;
        rom_memory[42131] = 3'b110;
        rom_memory[42132] = 3'b110;
        rom_memory[42133] = 3'b110;
        rom_memory[42134] = 3'b110;
        rom_memory[42135] = 3'b110;
        rom_memory[42136] = 3'b110;
        rom_memory[42137] = 3'b110;
        rom_memory[42138] = 3'b110;
        rom_memory[42139] = 3'b110;
        rom_memory[42140] = 3'b110;
        rom_memory[42141] = 3'b110;
        rom_memory[42142] = 3'b110;
        rom_memory[42143] = 3'b110;
        rom_memory[42144] = 3'b110;
        rom_memory[42145] = 3'b110;
        rom_memory[42146] = 3'b110;
        rom_memory[42147] = 3'b110;
        rom_memory[42148] = 3'b110;
        rom_memory[42149] = 3'b110;
        rom_memory[42150] = 3'b110;
        rom_memory[42151] = 3'b110;
        rom_memory[42152] = 3'b110;
        rom_memory[42153] = 3'b110;
        rom_memory[42154] = 3'b110;
        rom_memory[42155] = 3'b110;
        rom_memory[42156] = 3'b110;
        rom_memory[42157] = 3'b110;
        rom_memory[42158] = 3'b110;
        rom_memory[42159] = 3'b110;
        rom_memory[42160] = 3'b110;
        rom_memory[42161] = 3'b110;
        rom_memory[42162] = 3'b110;
        rom_memory[42163] = 3'b110;
        rom_memory[42164] = 3'b110;
        rom_memory[42165] = 3'b110;
        rom_memory[42166] = 3'b110;
        rom_memory[42167] = 3'b110;
        rom_memory[42168] = 3'b110;
        rom_memory[42169] = 3'b110;
        rom_memory[42170] = 3'b110;
        rom_memory[42171] = 3'b110;
        rom_memory[42172] = 3'b110;
        rom_memory[42173] = 3'b110;
        rom_memory[42174] = 3'b110;
        rom_memory[42175] = 3'b110;
        rom_memory[42176] = 3'b110;
        rom_memory[42177] = 3'b110;
        rom_memory[42178] = 3'b110;
        rom_memory[42179] = 3'b110;
        rom_memory[42180] = 3'b110;
        rom_memory[42181] = 3'b000;
        rom_memory[42182] = 3'b000;
        rom_memory[42183] = 3'b000;
        rom_memory[42184] = 3'b000;
        rom_memory[42185] = 3'b000;
        rom_memory[42186] = 3'b000;
        rom_memory[42187] = 3'b000;
        rom_memory[42188] = 3'b000;
        rom_memory[42189] = 3'b000;
        rom_memory[42190] = 3'b000;
        rom_memory[42191] = 3'b000;
        rom_memory[42192] = 3'b000;
        rom_memory[42193] = 3'b000;
        rom_memory[42194] = 3'b000;
        rom_memory[42195] = 3'b000;
        rom_memory[42196] = 3'b110;
        rom_memory[42197] = 3'b111;
        rom_memory[42198] = 3'b110;
        rom_memory[42199] = 3'b110;
        rom_memory[42200] = 3'b110;
        rom_memory[42201] = 3'b110;
        rom_memory[42202] = 3'b110;
        rom_memory[42203] = 3'b110;
        rom_memory[42204] = 3'b110;
        rom_memory[42205] = 3'b110;
        rom_memory[42206] = 3'b110;
        rom_memory[42207] = 3'b110;
        rom_memory[42208] = 3'b110;
        rom_memory[42209] = 3'b110;
        rom_memory[42210] = 3'b110;
        rom_memory[42211] = 3'b110;
        rom_memory[42212] = 3'b110;
        rom_memory[42213] = 3'b110;
        rom_memory[42214] = 3'b110;
        rom_memory[42215] = 3'b110;
        rom_memory[42216] = 3'b110;
        rom_memory[42217] = 3'b110;
        rom_memory[42218] = 3'b110;
        rom_memory[42219] = 3'b110;
        rom_memory[42220] = 3'b110;
        rom_memory[42221] = 3'b110;
        rom_memory[42222] = 3'b110;
        rom_memory[42223] = 3'b110;
        rom_memory[42224] = 3'b110;
        rom_memory[42225] = 3'b110;
        rom_memory[42226] = 3'b110;
        rom_memory[42227] = 3'b110;
        rom_memory[42228] = 3'b110;
        rom_memory[42229] = 3'b110;
        rom_memory[42230] = 3'b110;
        rom_memory[42231] = 3'b110;
        rom_memory[42232] = 3'b110;
        rom_memory[42233] = 3'b110;
        rom_memory[42234] = 3'b110;
        rom_memory[42235] = 3'b110;
        rom_memory[42236] = 3'b110;
        rom_memory[42237] = 3'b110;
        rom_memory[42238] = 3'b110;
        rom_memory[42239] = 3'b110;
        rom_memory[42240] = 3'b110;
        rom_memory[42241] = 3'b110;
        rom_memory[42242] = 3'b110;
        rom_memory[42243] = 3'b110;
        rom_memory[42244] = 3'b110;
        rom_memory[42245] = 3'b110;
        rom_memory[42246] = 3'b111;
        rom_memory[42247] = 3'b111;
        rom_memory[42248] = 3'b111;
        rom_memory[42249] = 3'b111;
        rom_memory[42250] = 3'b111;
        rom_memory[42251] = 3'b111;
        rom_memory[42252] = 3'b111;
        rom_memory[42253] = 3'b111;
        rom_memory[42254] = 3'b111;
        rom_memory[42255] = 3'b111;
        rom_memory[42256] = 3'b111;
        rom_memory[42257] = 3'b111;
        rom_memory[42258] = 3'b111;
        rom_memory[42259] = 3'b111;
        rom_memory[42260] = 3'b110;
        rom_memory[42261] = 3'b110;
        rom_memory[42262] = 3'b110;
        rom_memory[42263] = 3'b110;
        rom_memory[42264] = 3'b110;
        rom_memory[42265] = 3'b110;
        rom_memory[42266] = 3'b110;
        rom_memory[42267] = 3'b110;
        rom_memory[42268] = 3'b110;
        rom_memory[42269] = 3'b110;
        rom_memory[42270] = 3'b110;
        rom_memory[42271] = 3'b110;
        rom_memory[42272] = 3'b110;
        rom_memory[42273] = 3'b110;
        rom_memory[42274] = 3'b110;
        rom_memory[42275] = 3'b110;
        rom_memory[42276] = 3'b111;
        rom_memory[42277] = 3'b111;
        rom_memory[42278] = 3'b111;
        rom_memory[42279] = 3'b111;
        rom_memory[42280] = 3'b111;
        rom_memory[42281] = 3'b111;
        rom_memory[42282] = 3'b111;
        rom_memory[42283] = 3'b111;
        rom_memory[42284] = 3'b110;
        rom_memory[42285] = 3'b111;
        rom_memory[42286] = 3'b111;
        rom_memory[42287] = 3'b111;
        rom_memory[42288] = 3'b111;
        rom_memory[42289] = 3'b111;
        rom_memory[42290] = 3'b111;
        rom_memory[42291] = 3'b111;
        rom_memory[42292] = 3'b110;
        rom_memory[42293] = 3'b111;
        rom_memory[42294] = 3'b110;
        rom_memory[42295] = 3'b111;
        rom_memory[42296] = 3'b111;
        rom_memory[42297] = 3'b111;
        rom_memory[42298] = 3'b100;
        rom_memory[42299] = 3'b110;
        rom_memory[42300] = 3'b110;
        rom_memory[42301] = 3'b110;
        rom_memory[42302] = 3'b111;
        rom_memory[42303] = 3'b111;
        rom_memory[42304] = 3'b110;
        rom_memory[42305] = 3'b110;
        rom_memory[42306] = 3'b110;
        rom_memory[42307] = 3'b110;
        rom_memory[42308] = 3'b111;
        rom_memory[42309] = 3'b111;
        rom_memory[42310] = 3'b111;
        rom_memory[42311] = 3'b111;
        rom_memory[42312] = 3'b110;
        rom_memory[42313] = 3'b111;
        rom_memory[42314] = 3'b000;
        rom_memory[42315] = 3'b110;
        rom_memory[42316] = 3'b100;
        rom_memory[42317] = 3'b111;
        rom_memory[42318] = 3'b111;
        rom_memory[42319] = 3'b110;
        rom_memory[42320] = 3'b110;
        rom_memory[42321] = 3'b111;
        rom_memory[42322] = 3'b111;
        rom_memory[42323] = 3'b111;
        rom_memory[42324] = 3'b111;
        rom_memory[42325] = 3'b111;
        rom_memory[42326] = 3'b111;
        rom_memory[42327] = 3'b111;
        rom_memory[42328] = 3'b111;
        rom_memory[42329] = 3'b111;
        rom_memory[42330] = 3'b111;
        rom_memory[42331] = 3'b111;
        rom_memory[42332] = 3'b110;
        rom_memory[42333] = 3'b110;
        rom_memory[42334] = 3'b110;
        rom_memory[42335] = 3'b110;
        rom_memory[42336] = 3'b110;
        rom_memory[42337] = 3'b110;
        rom_memory[42338] = 3'b110;
        rom_memory[42339] = 3'b110;
        rom_memory[42340] = 3'b110;
        rom_memory[42341] = 3'b110;
        rom_memory[42342] = 3'b111;
        rom_memory[42343] = 3'b111;
        rom_memory[42344] = 3'b111;
        rom_memory[42345] = 3'b111;
        rom_memory[42346] = 3'b111;
        rom_memory[42347] = 3'b111;
        rom_memory[42348] = 3'b111;
        rom_memory[42349] = 3'b111;
        rom_memory[42350] = 3'b111;
        rom_memory[42351] = 3'b110;
        rom_memory[42352] = 3'b110;
        rom_memory[42353] = 3'b110;
        rom_memory[42354] = 3'b110;
        rom_memory[42355] = 3'b110;
        rom_memory[42356] = 3'b110;
        rom_memory[42357] = 3'b110;
        rom_memory[42358] = 3'b110;
        rom_memory[42359] = 3'b110;
        rom_memory[42360] = 3'b110;
        rom_memory[42361] = 3'b110;
        rom_memory[42362] = 3'b110;
        rom_memory[42363] = 3'b110;
        rom_memory[42364] = 3'b110;
        rom_memory[42365] = 3'b110;
        rom_memory[42366] = 3'b110;
        rom_memory[42367] = 3'b110;
        rom_memory[42368] = 3'b110;
        rom_memory[42369] = 3'b110;
        rom_memory[42370] = 3'b110;
        rom_memory[42371] = 3'b110;
        rom_memory[42372] = 3'b110;
        rom_memory[42373] = 3'b110;
        rom_memory[42374] = 3'b110;
        rom_memory[42375] = 3'b110;
        rom_memory[42376] = 3'b110;
        rom_memory[42377] = 3'b110;
        rom_memory[42378] = 3'b110;
        rom_memory[42379] = 3'b110;
        rom_memory[42380] = 3'b110;
        rom_memory[42381] = 3'b110;
        rom_memory[42382] = 3'b110;
        rom_memory[42383] = 3'b110;
        rom_memory[42384] = 3'b110;
        rom_memory[42385] = 3'b110;
        rom_memory[42386] = 3'b110;
        rom_memory[42387] = 3'b110;
        rom_memory[42388] = 3'b110;
        rom_memory[42389] = 3'b110;
        rom_memory[42390] = 3'b110;
        rom_memory[42391] = 3'b110;
        rom_memory[42392] = 3'b110;
        rom_memory[42393] = 3'b110;
        rom_memory[42394] = 3'b110;
        rom_memory[42395] = 3'b110;
        rom_memory[42396] = 3'b110;
        rom_memory[42397] = 3'b110;
        rom_memory[42398] = 3'b110;
        rom_memory[42399] = 3'b110;
        rom_memory[42400] = 3'b110;
        rom_memory[42401] = 3'b110;
        rom_memory[42402] = 3'b110;
        rom_memory[42403] = 3'b110;
        rom_memory[42404] = 3'b110;
        rom_memory[42405] = 3'b110;
        rom_memory[42406] = 3'b110;
        rom_memory[42407] = 3'b110;
        rom_memory[42408] = 3'b110;
        rom_memory[42409] = 3'b110;
        rom_memory[42410] = 3'b110;
        rom_memory[42411] = 3'b110;
        rom_memory[42412] = 3'b110;
        rom_memory[42413] = 3'b110;
        rom_memory[42414] = 3'b110;
        rom_memory[42415] = 3'b110;
        rom_memory[42416] = 3'b110;
        rom_memory[42417] = 3'b110;
        rom_memory[42418] = 3'b110;
        rom_memory[42419] = 3'b110;
        rom_memory[42420] = 3'b110;
        rom_memory[42421] = 3'b110;
        rom_memory[42422] = 3'b110;
        rom_memory[42423] = 3'b000;
        rom_memory[42424] = 3'b000;
        rom_memory[42425] = 3'b000;
        rom_memory[42426] = 3'b000;
        rom_memory[42427] = 3'b000;
        rom_memory[42428] = 3'b000;
        rom_memory[42429] = 3'b000;
        rom_memory[42430] = 3'b000;
        rom_memory[42431] = 3'b000;
        rom_memory[42432] = 3'b000;
        rom_memory[42433] = 3'b000;
        rom_memory[42434] = 3'b000;
        rom_memory[42435] = 3'b000;
        rom_memory[42436] = 3'b000;
        rom_memory[42437] = 3'b110;
        rom_memory[42438] = 3'b110;
        rom_memory[42439] = 3'b111;
        rom_memory[42440] = 3'b110;
        rom_memory[42441] = 3'b110;
        rom_memory[42442] = 3'b110;
        rom_memory[42443] = 3'b110;
        rom_memory[42444] = 3'b110;
        rom_memory[42445] = 3'b110;
        rom_memory[42446] = 3'b110;
        rom_memory[42447] = 3'b110;
        rom_memory[42448] = 3'b110;
        rom_memory[42449] = 3'b110;
        rom_memory[42450] = 3'b110;
        rom_memory[42451] = 3'b110;
        rom_memory[42452] = 3'b110;
        rom_memory[42453] = 3'b110;
        rom_memory[42454] = 3'b110;
        rom_memory[42455] = 3'b110;
        rom_memory[42456] = 3'b110;
        rom_memory[42457] = 3'b110;
        rom_memory[42458] = 3'b110;
        rom_memory[42459] = 3'b110;
        rom_memory[42460] = 3'b110;
        rom_memory[42461] = 3'b110;
        rom_memory[42462] = 3'b110;
        rom_memory[42463] = 3'b110;
        rom_memory[42464] = 3'b110;
        rom_memory[42465] = 3'b110;
        rom_memory[42466] = 3'b110;
        rom_memory[42467] = 3'b110;
        rom_memory[42468] = 3'b110;
        rom_memory[42469] = 3'b110;
        rom_memory[42470] = 3'b110;
        rom_memory[42471] = 3'b110;
        rom_memory[42472] = 3'b110;
        rom_memory[42473] = 3'b110;
        rom_memory[42474] = 3'b110;
        rom_memory[42475] = 3'b110;
        rom_memory[42476] = 3'b110;
        rom_memory[42477] = 3'b110;
        rom_memory[42478] = 3'b110;
        rom_memory[42479] = 3'b110;
        rom_memory[42480] = 3'b110;
        rom_memory[42481] = 3'b110;
        rom_memory[42482] = 3'b110;
        rom_memory[42483] = 3'b110;
        rom_memory[42484] = 3'b110;
        rom_memory[42485] = 3'b110;
        rom_memory[42486] = 3'b111;
        rom_memory[42487] = 3'b111;
        rom_memory[42488] = 3'b111;
        rom_memory[42489] = 3'b111;
        rom_memory[42490] = 3'b111;
        rom_memory[42491] = 3'b111;
        rom_memory[42492] = 3'b111;
        rom_memory[42493] = 3'b111;
        rom_memory[42494] = 3'b111;
        rom_memory[42495] = 3'b111;
        rom_memory[42496] = 3'b111;
        rom_memory[42497] = 3'b111;
        rom_memory[42498] = 3'b111;
        rom_memory[42499] = 3'b111;
        rom_memory[42500] = 3'b110;
        rom_memory[42501] = 3'b110;
        rom_memory[42502] = 3'b110;
        rom_memory[42503] = 3'b110;
        rom_memory[42504] = 3'b110;
        rom_memory[42505] = 3'b110;
        rom_memory[42506] = 3'b110;
        rom_memory[42507] = 3'b110;
        rom_memory[42508] = 3'b110;
        rom_memory[42509] = 3'b110;
        rom_memory[42510] = 3'b110;
        rom_memory[42511] = 3'b110;
        rom_memory[42512] = 3'b110;
        rom_memory[42513] = 3'b110;
        rom_memory[42514] = 3'b110;
        rom_memory[42515] = 3'b111;
        rom_memory[42516] = 3'b111;
        rom_memory[42517] = 3'b111;
        rom_memory[42518] = 3'b111;
        rom_memory[42519] = 3'b111;
        rom_memory[42520] = 3'b111;
        rom_memory[42521] = 3'b111;
        rom_memory[42522] = 3'b111;
        rom_memory[42523] = 3'b111;
        rom_memory[42524] = 3'b111;
        rom_memory[42525] = 3'b111;
        rom_memory[42526] = 3'b111;
        rom_memory[42527] = 3'b111;
        rom_memory[42528] = 3'b111;
        rom_memory[42529] = 3'b111;
        rom_memory[42530] = 3'b110;
        rom_memory[42531] = 3'b111;
        rom_memory[42532] = 3'b111;
        rom_memory[42533] = 3'b111;
        rom_memory[42534] = 3'b111;
        rom_memory[42535] = 3'b111;
        rom_memory[42536] = 3'b111;
        rom_memory[42537] = 3'b111;
        rom_memory[42538] = 3'b110;
        rom_memory[42539] = 3'b110;
        rom_memory[42540] = 3'b110;
        rom_memory[42541] = 3'b110;
        rom_memory[42542] = 3'b111;
        rom_memory[42543] = 3'b111;
        rom_memory[42544] = 3'b111;
        rom_memory[42545] = 3'b110;
        rom_memory[42546] = 3'b110;
        rom_memory[42547] = 3'b111;
        rom_memory[42548] = 3'b111;
        rom_memory[42549] = 3'b111;
        rom_memory[42550] = 3'b111;
        rom_memory[42551] = 3'b111;
        rom_memory[42552] = 3'b111;
        rom_memory[42553] = 3'b111;
        rom_memory[42554] = 3'b100;
        rom_memory[42555] = 3'b111;
        rom_memory[42556] = 3'b110;
        rom_memory[42557] = 3'b111;
        rom_memory[42558] = 3'b110;
        rom_memory[42559] = 3'b110;
        rom_memory[42560] = 3'b110;
        rom_memory[42561] = 3'b111;
        rom_memory[42562] = 3'b111;
        rom_memory[42563] = 3'b111;
        rom_memory[42564] = 3'b111;
        rom_memory[42565] = 3'b111;
        rom_memory[42566] = 3'b111;
        rom_memory[42567] = 3'b111;
        rom_memory[42568] = 3'b111;
        rom_memory[42569] = 3'b111;
        rom_memory[42570] = 3'b111;
        rom_memory[42571] = 3'b111;
        rom_memory[42572] = 3'b110;
        rom_memory[42573] = 3'b110;
        rom_memory[42574] = 3'b110;
        rom_memory[42575] = 3'b110;
        rom_memory[42576] = 3'b110;
        rom_memory[42577] = 3'b110;
        rom_memory[42578] = 3'b110;
        rom_memory[42579] = 3'b110;
        rom_memory[42580] = 3'b110;
        rom_memory[42581] = 3'b110;
        rom_memory[42582] = 3'b111;
        rom_memory[42583] = 3'b111;
        rom_memory[42584] = 3'b111;
        rom_memory[42585] = 3'b111;
        rom_memory[42586] = 3'b111;
        rom_memory[42587] = 3'b111;
        rom_memory[42588] = 3'b111;
        rom_memory[42589] = 3'b111;
        rom_memory[42590] = 3'b111;
        rom_memory[42591] = 3'b111;
        rom_memory[42592] = 3'b110;
        rom_memory[42593] = 3'b110;
        rom_memory[42594] = 3'b110;
        rom_memory[42595] = 3'b110;
        rom_memory[42596] = 3'b110;
        rom_memory[42597] = 3'b110;
        rom_memory[42598] = 3'b110;
        rom_memory[42599] = 3'b110;
        rom_memory[42600] = 3'b110;
        rom_memory[42601] = 3'b110;
        rom_memory[42602] = 3'b110;
        rom_memory[42603] = 3'b110;
        rom_memory[42604] = 3'b110;
        rom_memory[42605] = 3'b110;
        rom_memory[42606] = 3'b110;
        rom_memory[42607] = 3'b110;
        rom_memory[42608] = 3'b110;
        rom_memory[42609] = 3'b110;
        rom_memory[42610] = 3'b110;
        rom_memory[42611] = 3'b110;
        rom_memory[42612] = 3'b110;
        rom_memory[42613] = 3'b110;
        rom_memory[42614] = 3'b110;
        rom_memory[42615] = 3'b110;
        rom_memory[42616] = 3'b110;
        rom_memory[42617] = 3'b110;
        rom_memory[42618] = 3'b110;
        rom_memory[42619] = 3'b110;
        rom_memory[42620] = 3'b110;
        rom_memory[42621] = 3'b110;
        rom_memory[42622] = 3'b110;
        rom_memory[42623] = 3'b110;
        rom_memory[42624] = 3'b110;
        rom_memory[42625] = 3'b110;
        rom_memory[42626] = 3'b110;
        rom_memory[42627] = 3'b110;
        rom_memory[42628] = 3'b110;
        rom_memory[42629] = 3'b110;
        rom_memory[42630] = 3'b110;
        rom_memory[42631] = 3'b110;
        rom_memory[42632] = 3'b110;
        rom_memory[42633] = 3'b110;
        rom_memory[42634] = 3'b110;
        rom_memory[42635] = 3'b110;
        rom_memory[42636] = 3'b110;
        rom_memory[42637] = 3'b110;
        rom_memory[42638] = 3'b110;
        rom_memory[42639] = 3'b110;
        rom_memory[42640] = 3'b110;
        rom_memory[42641] = 3'b110;
        rom_memory[42642] = 3'b110;
        rom_memory[42643] = 3'b110;
        rom_memory[42644] = 3'b110;
        rom_memory[42645] = 3'b110;
        rom_memory[42646] = 3'b110;
        rom_memory[42647] = 3'b110;
        rom_memory[42648] = 3'b110;
        rom_memory[42649] = 3'b110;
        rom_memory[42650] = 3'b110;
        rom_memory[42651] = 3'b110;
        rom_memory[42652] = 3'b110;
        rom_memory[42653] = 3'b110;
        rom_memory[42654] = 3'b110;
        rom_memory[42655] = 3'b110;
        rom_memory[42656] = 3'b110;
        rom_memory[42657] = 3'b110;
        rom_memory[42658] = 3'b110;
        rom_memory[42659] = 3'b110;
        rom_memory[42660] = 3'b110;
        rom_memory[42661] = 3'b110;
        rom_memory[42662] = 3'b110;
        rom_memory[42663] = 3'b110;
        rom_memory[42664] = 3'b110;
        rom_memory[42665] = 3'b000;
        rom_memory[42666] = 3'b000;
        rom_memory[42667] = 3'b000;
        rom_memory[42668] = 3'b000;
        rom_memory[42669] = 3'b000;
        rom_memory[42670] = 3'b000;
        rom_memory[42671] = 3'b000;
        rom_memory[42672] = 3'b000;
        rom_memory[42673] = 3'b000;
        rom_memory[42674] = 3'b000;
        rom_memory[42675] = 3'b000;
        rom_memory[42676] = 3'b000;
        rom_memory[42677] = 3'b000;
        rom_memory[42678] = 3'b000;
        rom_memory[42679] = 3'b110;
        rom_memory[42680] = 3'b110;
        rom_memory[42681] = 3'b110;
        rom_memory[42682] = 3'b110;
        rom_memory[42683] = 3'b110;
        rom_memory[42684] = 3'b110;
        rom_memory[42685] = 3'b110;
        rom_memory[42686] = 3'b110;
        rom_memory[42687] = 3'b110;
        rom_memory[42688] = 3'b110;
        rom_memory[42689] = 3'b110;
        rom_memory[42690] = 3'b110;
        rom_memory[42691] = 3'b110;
        rom_memory[42692] = 3'b110;
        rom_memory[42693] = 3'b110;
        rom_memory[42694] = 3'b110;
        rom_memory[42695] = 3'b110;
        rom_memory[42696] = 3'b110;
        rom_memory[42697] = 3'b110;
        rom_memory[42698] = 3'b110;
        rom_memory[42699] = 3'b110;
        rom_memory[42700] = 3'b110;
        rom_memory[42701] = 3'b110;
        rom_memory[42702] = 3'b110;
        rom_memory[42703] = 3'b110;
        rom_memory[42704] = 3'b110;
        rom_memory[42705] = 3'b110;
        rom_memory[42706] = 3'b110;
        rom_memory[42707] = 3'b110;
        rom_memory[42708] = 3'b110;
        rom_memory[42709] = 3'b110;
        rom_memory[42710] = 3'b110;
        rom_memory[42711] = 3'b110;
        rom_memory[42712] = 3'b110;
        rom_memory[42713] = 3'b110;
        rom_memory[42714] = 3'b110;
        rom_memory[42715] = 3'b110;
        rom_memory[42716] = 3'b110;
        rom_memory[42717] = 3'b110;
        rom_memory[42718] = 3'b110;
        rom_memory[42719] = 3'b110;
        rom_memory[42720] = 3'b110;
        rom_memory[42721] = 3'b110;
        rom_memory[42722] = 3'b110;
        rom_memory[42723] = 3'b110;
        rom_memory[42724] = 3'b111;
        rom_memory[42725] = 3'b111;
        rom_memory[42726] = 3'b111;
        rom_memory[42727] = 3'b111;
        rom_memory[42728] = 3'b111;
        rom_memory[42729] = 3'b111;
        rom_memory[42730] = 3'b111;
        rom_memory[42731] = 3'b111;
        rom_memory[42732] = 3'b111;
        rom_memory[42733] = 3'b111;
        rom_memory[42734] = 3'b111;
        rom_memory[42735] = 3'b111;
        rom_memory[42736] = 3'b111;
        rom_memory[42737] = 3'b111;
        rom_memory[42738] = 3'b111;
        rom_memory[42739] = 3'b111;
        rom_memory[42740] = 3'b110;
        rom_memory[42741] = 3'b110;
        rom_memory[42742] = 3'b110;
        rom_memory[42743] = 3'b110;
        rom_memory[42744] = 3'b110;
        rom_memory[42745] = 3'b110;
        rom_memory[42746] = 3'b110;
        rom_memory[42747] = 3'b110;
        rom_memory[42748] = 3'b110;
        rom_memory[42749] = 3'b110;
        rom_memory[42750] = 3'b110;
        rom_memory[42751] = 3'b110;
        rom_memory[42752] = 3'b110;
        rom_memory[42753] = 3'b110;
        rom_memory[42754] = 3'b111;
        rom_memory[42755] = 3'b111;
        rom_memory[42756] = 3'b111;
        rom_memory[42757] = 3'b111;
        rom_memory[42758] = 3'b111;
        rom_memory[42759] = 3'b111;
        rom_memory[42760] = 3'b111;
        rom_memory[42761] = 3'b111;
        rom_memory[42762] = 3'b111;
        rom_memory[42763] = 3'b111;
        rom_memory[42764] = 3'b111;
        rom_memory[42765] = 3'b111;
        rom_memory[42766] = 3'b111;
        rom_memory[42767] = 3'b111;
        rom_memory[42768] = 3'b111;
        rom_memory[42769] = 3'b111;
        rom_memory[42770] = 3'b111;
        rom_memory[42771] = 3'b111;
        rom_memory[42772] = 3'b111;
        rom_memory[42773] = 3'b111;
        rom_memory[42774] = 3'b111;
        rom_memory[42775] = 3'b111;
        rom_memory[42776] = 3'b111;
        rom_memory[42777] = 3'b111;
        rom_memory[42778] = 3'b110;
        rom_memory[42779] = 3'b110;
        rom_memory[42780] = 3'b110;
        rom_memory[42781] = 3'b110;
        rom_memory[42782] = 3'b111;
        rom_memory[42783] = 3'b110;
        rom_memory[42784] = 3'b111;
        rom_memory[42785] = 3'b111;
        rom_memory[42786] = 3'b111;
        rom_memory[42787] = 3'b111;
        rom_memory[42788] = 3'b110;
        rom_memory[42789] = 3'b110;
        rom_memory[42790] = 3'b110;
        rom_memory[42791] = 3'b111;
        rom_memory[42792] = 3'b111;
        rom_memory[42793] = 3'b111;
        rom_memory[42794] = 3'b000;
        rom_memory[42795] = 3'b111;
        rom_memory[42796] = 3'b110;
        rom_memory[42797] = 3'b110;
        rom_memory[42798] = 3'b110;
        rom_memory[42799] = 3'b110;
        rom_memory[42800] = 3'b111;
        rom_memory[42801] = 3'b110;
        rom_memory[42802] = 3'b111;
        rom_memory[42803] = 3'b110;
        rom_memory[42804] = 3'b100;
        rom_memory[42805] = 3'b111;
        rom_memory[42806] = 3'b111;
        rom_memory[42807] = 3'b111;
        rom_memory[42808] = 3'b111;
        rom_memory[42809] = 3'b111;
        rom_memory[42810] = 3'b110;
        rom_memory[42811] = 3'b110;
        rom_memory[42812] = 3'b110;
        rom_memory[42813] = 3'b111;
        rom_memory[42814] = 3'b111;
        rom_memory[42815] = 3'b111;
        rom_memory[42816] = 3'b110;
        rom_memory[42817] = 3'b110;
        rom_memory[42818] = 3'b110;
        rom_memory[42819] = 3'b110;
        rom_memory[42820] = 3'b110;
        rom_memory[42821] = 3'b110;
        rom_memory[42822] = 3'b110;
        rom_memory[42823] = 3'b111;
        rom_memory[42824] = 3'b111;
        rom_memory[42825] = 3'b111;
        rom_memory[42826] = 3'b111;
        rom_memory[42827] = 3'b111;
        rom_memory[42828] = 3'b111;
        rom_memory[42829] = 3'b111;
        rom_memory[42830] = 3'b111;
        rom_memory[42831] = 3'b111;
        rom_memory[42832] = 3'b110;
        rom_memory[42833] = 3'b110;
        rom_memory[42834] = 3'b110;
        rom_memory[42835] = 3'b110;
        rom_memory[42836] = 3'b110;
        rom_memory[42837] = 3'b110;
        rom_memory[42838] = 3'b110;
        rom_memory[42839] = 3'b110;
        rom_memory[42840] = 3'b110;
        rom_memory[42841] = 3'b110;
        rom_memory[42842] = 3'b110;
        rom_memory[42843] = 3'b110;
        rom_memory[42844] = 3'b110;
        rom_memory[42845] = 3'b110;
        rom_memory[42846] = 3'b110;
        rom_memory[42847] = 3'b110;
        rom_memory[42848] = 3'b110;
        rom_memory[42849] = 3'b110;
        rom_memory[42850] = 3'b110;
        rom_memory[42851] = 3'b110;
        rom_memory[42852] = 3'b110;
        rom_memory[42853] = 3'b110;
        rom_memory[42854] = 3'b110;
        rom_memory[42855] = 3'b110;
        rom_memory[42856] = 3'b110;
        rom_memory[42857] = 3'b110;
        rom_memory[42858] = 3'b110;
        rom_memory[42859] = 3'b110;
        rom_memory[42860] = 3'b110;
        rom_memory[42861] = 3'b110;
        rom_memory[42862] = 3'b110;
        rom_memory[42863] = 3'b110;
        rom_memory[42864] = 3'b110;
        rom_memory[42865] = 3'b110;
        rom_memory[42866] = 3'b110;
        rom_memory[42867] = 3'b110;
        rom_memory[42868] = 3'b110;
        rom_memory[42869] = 3'b110;
        rom_memory[42870] = 3'b110;
        rom_memory[42871] = 3'b110;
        rom_memory[42872] = 3'b110;
        rom_memory[42873] = 3'b110;
        rom_memory[42874] = 3'b110;
        rom_memory[42875] = 3'b110;
        rom_memory[42876] = 3'b110;
        rom_memory[42877] = 3'b110;
        rom_memory[42878] = 3'b110;
        rom_memory[42879] = 3'b110;
        rom_memory[42880] = 3'b110;
        rom_memory[42881] = 3'b110;
        rom_memory[42882] = 3'b110;
        rom_memory[42883] = 3'b110;
        rom_memory[42884] = 3'b110;
        rom_memory[42885] = 3'b110;
        rom_memory[42886] = 3'b110;
        rom_memory[42887] = 3'b110;
        rom_memory[42888] = 3'b110;
        rom_memory[42889] = 3'b110;
        rom_memory[42890] = 3'b110;
        rom_memory[42891] = 3'b110;
        rom_memory[42892] = 3'b110;
        rom_memory[42893] = 3'b110;
        rom_memory[42894] = 3'b110;
        rom_memory[42895] = 3'b110;
        rom_memory[42896] = 3'b110;
        rom_memory[42897] = 3'b110;
        rom_memory[42898] = 3'b110;
        rom_memory[42899] = 3'b110;
        rom_memory[42900] = 3'b110;
        rom_memory[42901] = 3'b110;
        rom_memory[42902] = 3'b110;
        rom_memory[42903] = 3'b110;
        rom_memory[42904] = 3'b110;
        rom_memory[42905] = 3'b110;
        rom_memory[42906] = 3'b110;
        rom_memory[42907] = 3'b000;
        rom_memory[42908] = 3'b000;
        rom_memory[42909] = 3'b000;
        rom_memory[42910] = 3'b000;
        rom_memory[42911] = 3'b000;
        rom_memory[42912] = 3'b000;
        rom_memory[42913] = 3'b000;
        rom_memory[42914] = 3'b000;
        rom_memory[42915] = 3'b000;
        rom_memory[42916] = 3'b000;
        rom_memory[42917] = 3'b000;
        rom_memory[42918] = 3'b000;
        rom_memory[42919] = 3'b000;
        rom_memory[42920] = 3'b100;
        rom_memory[42921] = 3'b111;
        rom_memory[42922] = 3'b111;
        rom_memory[42923] = 3'b110;
        rom_memory[42924] = 3'b110;
        rom_memory[42925] = 3'b110;
        rom_memory[42926] = 3'b110;
        rom_memory[42927] = 3'b110;
        rom_memory[42928] = 3'b110;
        rom_memory[42929] = 3'b110;
        rom_memory[42930] = 3'b110;
        rom_memory[42931] = 3'b110;
        rom_memory[42932] = 3'b110;
        rom_memory[42933] = 3'b110;
        rom_memory[42934] = 3'b110;
        rom_memory[42935] = 3'b110;
        rom_memory[42936] = 3'b110;
        rom_memory[42937] = 3'b110;
        rom_memory[42938] = 3'b110;
        rom_memory[42939] = 3'b110;
        rom_memory[42940] = 3'b110;
        rom_memory[42941] = 3'b110;
        rom_memory[42942] = 3'b110;
        rom_memory[42943] = 3'b110;
        rom_memory[42944] = 3'b110;
        rom_memory[42945] = 3'b110;
        rom_memory[42946] = 3'b110;
        rom_memory[42947] = 3'b110;
        rom_memory[42948] = 3'b110;
        rom_memory[42949] = 3'b110;
        rom_memory[42950] = 3'b110;
        rom_memory[42951] = 3'b110;
        rom_memory[42952] = 3'b110;
        rom_memory[42953] = 3'b110;
        rom_memory[42954] = 3'b110;
        rom_memory[42955] = 3'b110;
        rom_memory[42956] = 3'b110;
        rom_memory[42957] = 3'b110;
        rom_memory[42958] = 3'b110;
        rom_memory[42959] = 3'b110;
        rom_memory[42960] = 3'b111;
        rom_memory[42961] = 3'b111;
        rom_memory[42962] = 3'b111;
        rom_memory[42963] = 3'b111;
        rom_memory[42964] = 3'b111;
        rom_memory[42965] = 3'b111;
        rom_memory[42966] = 3'b111;
        rom_memory[42967] = 3'b111;
        rom_memory[42968] = 3'b111;
        rom_memory[42969] = 3'b111;
        rom_memory[42970] = 3'b111;
        rom_memory[42971] = 3'b111;
        rom_memory[42972] = 3'b111;
        rom_memory[42973] = 3'b111;
        rom_memory[42974] = 3'b111;
        rom_memory[42975] = 3'b111;
        rom_memory[42976] = 3'b111;
        rom_memory[42977] = 3'b111;
        rom_memory[42978] = 3'b111;
        rom_memory[42979] = 3'b111;
        rom_memory[42980] = 3'b111;
        rom_memory[42981] = 3'b110;
        rom_memory[42982] = 3'b110;
        rom_memory[42983] = 3'b110;
        rom_memory[42984] = 3'b110;
        rom_memory[42985] = 3'b110;
        rom_memory[42986] = 3'b110;
        rom_memory[42987] = 3'b110;
        rom_memory[42988] = 3'b110;
        rom_memory[42989] = 3'b110;
        rom_memory[42990] = 3'b110;
        rom_memory[42991] = 3'b110;
        rom_memory[42992] = 3'b110;
        rom_memory[42993] = 3'b110;
        rom_memory[42994] = 3'b111;
        rom_memory[42995] = 3'b111;
        rom_memory[42996] = 3'b111;
        rom_memory[42997] = 3'b111;
        rom_memory[42998] = 3'b111;
        rom_memory[42999] = 3'b111;
        rom_memory[43000] = 3'b111;
        rom_memory[43001] = 3'b111;
        rom_memory[43002] = 3'b111;
        rom_memory[43003] = 3'b111;
        rom_memory[43004] = 3'b110;
        rom_memory[43005] = 3'b110;
        rom_memory[43006] = 3'b111;
        rom_memory[43007] = 3'b111;
        rom_memory[43008] = 3'b111;
        rom_memory[43009] = 3'b111;
        rom_memory[43010] = 3'b111;
        rom_memory[43011] = 3'b111;
        rom_memory[43012] = 3'b111;
        rom_memory[43013] = 3'b111;
        rom_memory[43014] = 3'b111;
        rom_memory[43015] = 3'b111;
        rom_memory[43016] = 3'b111;
        rom_memory[43017] = 3'b111;
        rom_memory[43018] = 3'b110;
        rom_memory[43019] = 3'b110;
        rom_memory[43020] = 3'b110;
        rom_memory[43021] = 3'b100;
        rom_memory[43022] = 3'b111;
        rom_memory[43023] = 3'b110;
        rom_memory[43024] = 3'b110;
        rom_memory[43025] = 3'b110;
        rom_memory[43026] = 3'b110;
        rom_memory[43027] = 3'b111;
        rom_memory[43028] = 3'b110;
        rom_memory[43029] = 3'b110;
        rom_memory[43030] = 3'b110;
        rom_memory[43031] = 3'b111;
        rom_memory[43032] = 3'b111;
        rom_memory[43033] = 3'b111;
        rom_memory[43034] = 3'b000;
        rom_memory[43035] = 3'b100;
        rom_memory[43036] = 3'b110;
        rom_memory[43037] = 3'b110;
        rom_memory[43038] = 3'b110;
        rom_memory[43039] = 3'b110;
        rom_memory[43040] = 3'b110;
        rom_memory[43041] = 3'b110;
        rom_memory[43042] = 3'b111;
        rom_memory[43043] = 3'b110;
        rom_memory[43044] = 3'b110;
        rom_memory[43045] = 3'b110;
        rom_memory[43046] = 3'b110;
        rom_memory[43047] = 3'b110;
        rom_memory[43048] = 3'b110;
        rom_memory[43049] = 3'b110;
        rom_memory[43050] = 3'b110;
        rom_memory[43051] = 3'b110;
        rom_memory[43052] = 3'b110;
        rom_memory[43053] = 3'b111;
        rom_memory[43054] = 3'b111;
        rom_memory[43055] = 3'b111;
        rom_memory[43056] = 3'b111;
        rom_memory[43057] = 3'b111;
        rom_memory[43058] = 3'b110;
        rom_memory[43059] = 3'b110;
        rom_memory[43060] = 3'b110;
        rom_memory[43061] = 3'b110;
        rom_memory[43062] = 3'b110;
        rom_memory[43063] = 3'b111;
        rom_memory[43064] = 3'b111;
        rom_memory[43065] = 3'b111;
        rom_memory[43066] = 3'b111;
        rom_memory[43067] = 3'b111;
        rom_memory[43068] = 3'b111;
        rom_memory[43069] = 3'b111;
        rom_memory[43070] = 3'b111;
        rom_memory[43071] = 3'b111;
        rom_memory[43072] = 3'b111;
        rom_memory[43073] = 3'b110;
        rom_memory[43074] = 3'b110;
        rom_memory[43075] = 3'b110;
        rom_memory[43076] = 3'b110;
        rom_memory[43077] = 3'b110;
        rom_memory[43078] = 3'b110;
        rom_memory[43079] = 3'b110;
        rom_memory[43080] = 3'b110;
        rom_memory[43081] = 3'b110;
        rom_memory[43082] = 3'b110;
        rom_memory[43083] = 3'b110;
        rom_memory[43084] = 3'b110;
        rom_memory[43085] = 3'b110;
        rom_memory[43086] = 3'b110;
        rom_memory[43087] = 3'b110;
        rom_memory[43088] = 3'b110;
        rom_memory[43089] = 3'b110;
        rom_memory[43090] = 3'b110;
        rom_memory[43091] = 3'b110;
        rom_memory[43092] = 3'b110;
        rom_memory[43093] = 3'b110;
        rom_memory[43094] = 3'b110;
        rom_memory[43095] = 3'b110;
        rom_memory[43096] = 3'b110;
        rom_memory[43097] = 3'b110;
        rom_memory[43098] = 3'b110;
        rom_memory[43099] = 3'b110;
        rom_memory[43100] = 3'b110;
        rom_memory[43101] = 3'b110;
        rom_memory[43102] = 3'b110;
        rom_memory[43103] = 3'b110;
        rom_memory[43104] = 3'b110;
        rom_memory[43105] = 3'b110;
        rom_memory[43106] = 3'b110;
        rom_memory[43107] = 3'b110;
        rom_memory[43108] = 3'b110;
        rom_memory[43109] = 3'b110;
        rom_memory[43110] = 3'b110;
        rom_memory[43111] = 3'b110;
        rom_memory[43112] = 3'b110;
        rom_memory[43113] = 3'b110;
        rom_memory[43114] = 3'b110;
        rom_memory[43115] = 3'b110;
        rom_memory[43116] = 3'b110;
        rom_memory[43117] = 3'b110;
        rom_memory[43118] = 3'b110;
        rom_memory[43119] = 3'b110;
        rom_memory[43120] = 3'b110;
        rom_memory[43121] = 3'b110;
        rom_memory[43122] = 3'b110;
        rom_memory[43123] = 3'b110;
        rom_memory[43124] = 3'b110;
        rom_memory[43125] = 3'b110;
        rom_memory[43126] = 3'b110;
        rom_memory[43127] = 3'b110;
        rom_memory[43128] = 3'b110;
        rom_memory[43129] = 3'b110;
        rom_memory[43130] = 3'b110;
        rom_memory[43131] = 3'b110;
        rom_memory[43132] = 3'b110;
        rom_memory[43133] = 3'b110;
        rom_memory[43134] = 3'b110;
        rom_memory[43135] = 3'b110;
        rom_memory[43136] = 3'b110;
        rom_memory[43137] = 3'b110;
        rom_memory[43138] = 3'b110;
        rom_memory[43139] = 3'b110;
        rom_memory[43140] = 3'b110;
        rom_memory[43141] = 3'b110;
        rom_memory[43142] = 3'b110;
        rom_memory[43143] = 3'b110;
        rom_memory[43144] = 3'b110;
        rom_memory[43145] = 3'b110;
        rom_memory[43146] = 3'b110;
        rom_memory[43147] = 3'b110;
        rom_memory[43148] = 3'b110;
        rom_memory[43149] = 3'b000;
        rom_memory[43150] = 3'b000;
        rom_memory[43151] = 3'b000;
        rom_memory[43152] = 3'b000;
        rom_memory[43153] = 3'b000;
        rom_memory[43154] = 3'b000;
        rom_memory[43155] = 3'b000;
        rom_memory[43156] = 3'b000;
        rom_memory[43157] = 3'b000;
        rom_memory[43158] = 3'b000;
        rom_memory[43159] = 3'b000;
        rom_memory[43160] = 3'b000;
        rom_memory[43161] = 3'b000;
        rom_memory[43162] = 3'b100;
        rom_memory[43163] = 3'b110;
        rom_memory[43164] = 3'b111;
        rom_memory[43165] = 3'b110;
        rom_memory[43166] = 3'b110;
        rom_memory[43167] = 3'b110;
        rom_memory[43168] = 3'b110;
        rom_memory[43169] = 3'b110;
        rom_memory[43170] = 3'b110;
        rom_memory[43171] = 3'b110;
        rom_memory[43172] = 3'b110;
        rom_memory[43173] = 3'b110;
        rom_memory[43174] = 3'b110;
        rom_memory[43175] = 3'b110;
        rom_memory[43176] = 3'b110;
        rom_memory[43177] = 3'b110;
        rom_memory[43178] = 3'b110;
        rom_memory[43179] = 3'b110;
        rom_memory[43180] = 3'b110;
        rom_memory[43181] = 3'b110;
        rom_memory[43182] = 3'b110;
        rom_memory[43183] = 3'b110;
        rom_memory[43184] = 3'b110;
        rom_memory[43185] = 3'b110;
        rom_memory[43186] = 3'b110;
        rom_memory[43187] = 3'b110;
        rom_memory[43188] = 3'b110;
        rom_memory[43189] = 3'b110;
        rom_memory[43190] = 3'b110;
        rom_memory[43191] = 3'b110;
        rom_memory[43192] = 3'b110;
        rom_memory[43193] = 3'b110;
        rom_memory[43194] = 3'b110;
        rom_memory[43195] = 3'b110;
        rom_memory[43196] = 3'b110;
        rom_memory[43197] = 3'b110;
        rom_memory[43198] = 3'b110;
        rom_memory[43199] = 3'b110;
        rom_memory[43200] = 3'b111;
        rom_memory[43201] = 3'b111;
        rom_memory[43202] = 3'b111;
        rom_memory[43203] = 3'b111;
        rom_memory[43204] = 3'b111;
        rom_memory[43205] = 3'b111;
        rom_memory[43206] = 3'b111;
        rom_memory[43207] = 3'b111;
        rom_memory[43208] = 3'b111;
        rom_memory[43209] = 3'b111;
        rom_memory[43210] = 3'b111;
        rom_memory[43211] = 3'b111;
        rom_memory[43212] = 3'b111;
        rom_memory[43213] = 3'b111;
        rom_memory[43214] = 3'b111;
        rom_memory[43215] = 3'b111;
        rom_memory[43216] = 3'b111;
        rom_memory[43217] = 3'b111;
        rom_memory[43218] = 3'b111;
        rom_memory[43219] = 3'b111;
        rom_memory[43220] = 3'b111;
        rom_memory[43221] = 3'b110;
        rom_memory[43222] = 3'b110;
        rom_memory[43223] = 3'b110;
        rom_memory[43224] = 3'b110;
        rom_memory[43225] = 3'b110;
        rom_memory[43226] = 3'b110;
        rom_memory[43227] = 3'b110;
        rom_memory[43228] = 3'b110;
        rom_memory[43229] = 3'b110;
        rom_memory[43230] = 3'b110;
        rom_memory[43231] = 3'b110;
        rom_memory[43232] = 3'b110;
        rom_memory[43233] = 3'b111;
        rom_memory[43234] = 3'b111;
        rom_memory[43235] = 3'b111;
        rom_memory[43236] = 3'b111;
        rom_memory[43237] = 3'b111;
        rom_memory[43238] = 3'b111;
        rom_memory[43239] = 3'b111;
        rom_memory[43240] = 3'b111;
        rom_memory[43241] = 3'b111;
        rom_memory[43242] = 3'b111;
        rom_memory[43243] = 3'b111;
        rom_memory[43244] = 3'b110;
        rom_memory[43245] = 3'b110;
        rom_memory[43246] = 3'b110;
        rom_memory[43247] = 3'b110;
        rom_memory[43248] = 3'b111;
        rom_memory[43249] = 3'b111;
        rom_memory[43250] = 3'b111;
        rom_memory[43251] = 3'b111;
        rom_memory[43252] = 3'b111;
        rom_memory[43253] = 3'b111;
        rom_memory[43254] = 3'b111;
        rom_memory[43255] = 3'b111;
        rom_memory[43256] = 3'b111;
        rom_memory[43257] = 3'b110;
        rom_memory[43258] = 3'b111;
        rom_memory[43259] = 3'b111;
        rom_memory[43260] = 3'b110;
        rom_memory[43261] = 3'b100;
        rom_memory[43262] = 3'b110;
        rom_memory[43263] = 3'b111;
        rom_memory[43264] = 3'b110;
        rom_memory[43265] = 3'b110;
        rom_memory[43266] = 3'b110;
        rom_memory[43267] = 3'b111;
        rom_memory[43268] = 3'b110;
        rom_memory[43269] = 3'b110;
        rom_memory[43270] = 3'b110;
        rom_memory[43271] = 3'b111;
        rom_memory[43272] = 3'b111;
        rom_memory[43273] = 3'b111;
        rom_memory[43274] = 3'b100;
        rom_memory[43275] = 3'b111;
        rom_memory[43276] = 3'b110;
        rom_memory[43277] = 3'b110;
        rom_memory[43278] = 3'b110;
        rom_memory[43279] = 3'b110;
        rom_memory[43280] = 3'b110;
        rom_memory[43281] = 3'b110;
        rom_memory[43282] = 3'b110;
        rom_memory[43283] = 3'b110;
        rom_memory[43284] = 3'b110;
        rom_memory[43285] = 3'b110;
        rom_memory[43286] = 3'b110;
        rom_memory[43287] = 3'b110;
        rom_memory[43288] = 3'b110;
        rom_memory[43289] = 3'b110;
        rom_memory[43290] = 3'b110;
        rom_memory[43291] = 3'b110;
        rom_memory[43292] = 3'b110;
        rom_memory[43293] = 3'b111;
        rom_memory[43294] = 3'b111;
        rom_memory[43295] = 3'b111;
        rom_memory[43296] = 3'b111;
        rom_memory[43297] = 3'b111;
        rom_memory[43298] = 3'b110;
        rom_memory[43299] = 3'b110;
        rom_memory[43300] = 3'b110;
        rom_memory[43301] = 3'b110;
        rom_memory[43302] = 3'b110;
        rom_memory[43303] = 3'b111;
        rom_memory[43304] = 3'b111;
        rom_memory[43305] = 3'b111;
        rom_memory[43306] = 3'b111;
        rom_memory[43307] = 3'b111;
        rom_memory[43308] = 3'b111;
        rom_memory[43309] = 3'b111;
        rom_memory[43310] = 3'b111;
        rom_memory[43311] = 3'b111;
        rom_memory[43312] = 3'b111;
        rom_memory[43313] = 3'b110;
        rom_memory[43314] = 3'b110;
        rom_memory[43315] = 3'b110;
        rom_memory[43316] = 3'b110;
        rom_memory[43317] = 3'b110;
        rom_memory[43318] = 3'b110;
        rom_memory[43319] = 3'b110;
        rom_memory[43320] = 3'b110;
        rom_memory[43321] = 3'b110;
        rom_memory[43322] = 3'b110;
        rom_memory[43323] = 3'b110;
        rom_memory[43324] = 3'b110;
        rom_memory[43325] = 3'b110;
        rom_memory[43326] = 3'b110;
        rom_memory[43327] = 3'b110;
        rom_memory[43328] = 3'b110;
        rom_memory[43329] = 3'b110;
        rom_memory[43330] = 3'b110;
        rom_memory[43331] = 3'b110;
        rom_memory[43332] = 3'b110;
        rom_memory[43333] = 3'b110;
        rom_memory[43334] = 3'b110;
        rom_memory[43335] = 3'b110;
        rom_memory[43336] = 3'b110;
        rom_memory[43337] = 3'b110;
        rom_memory[43338] = 3'b110;
        rom_memory[43339] = 3'b110;
        rom_memory[43340] = 3'b110;
        rom_memory[43341] = 3'b110;
        rom_memory[43342] = 3'b110;
        rom_memory[43343] = 3'b110;
        rom_memory[43344] = 3'b110;
        rom_memory[43345] = 3'b110;
        rom_memory[43346] = 3'b110;
        rom_memory[43347] = 3'b110;
        rom_memory[43348] = 3'b110;
        rom_memory[43349] = 3'b110;
        rom_memory[43350] = 3'b110;
        rom_memory[43351] = 3'b110;
        rom_memory[43352] = 3'b110;
        rom_memory[43353] = 3'b110;
        rom_memory[43354] = 3'b110;
        rom_memory[43355] = 3'b110;
        rom_memory[43356] = 3'b110;
        rom_memory[43357] = 3'b110;
        rom_memory[43358] = 3'b110;
        rom_memory[43359] = 3'b110;
        rom_memory[43360] = 3'b110;
        rom_memory[43361] = 3'b110;
        rom_memory[43362] = 3'b110;
        rom_memory[43363] = 3'b110;
        rom_memory[43364] = 3'b110;
        rom_memory[43365] = 3'b110;
        rom_memory[43366] = 3'b110;
        rom_memory[43367] = 3'b110;
        rom_memory[43368] = 3'b110;
        rom_memory[43369] = 3'b110;
        rom_memory[43370] = 3'b110;
        rom_memory[43371] = 3'b110;
        rom_memory[43372] = 3'b110;
        rom_memory[43373] = 3'b110;
        rom_memory[43374] = 3'b110;
        rom_memory[43375] = 3'b110;
        rom_memory[43376] = 3'b110;
        rom_memory[43377] = 3'b110;
        rom_memory[43378] = 3'b110;
        rom_memory[43379] = 3'b110;
        rom_memory[43380] = 3'b110;
        rom_memory[43381] = 3'b110;
        rom_memory[43382] = 3'b110;
        rom_memory[43383] = 3'b110;
        rom_memory[43384] = 3'b110;
        rom_memory[43385] = 3'b110;
        rom_memory[43386] = 3'b110;
        rom_memory[43387] = 3'b110;
        rom_memory[43388] = 3'b110;
        rom_memory[43389] = 3'b110;
        rom_memory[43390] = 3'b110;
        rom_memory[43391] = 3'b000;
        rom_memory[43392] = 3'b000;
        rom_memory[43393] = 3'b000;
        rom_memory[43394] = 3'b000;
        rom_memory[43395] = 3'b000;
        rom_memory[43396] = 3'b000;
        rom_memory[43397] = 3'b000;
        rom_memory[43398] = 3'b000;
        rom_memory[43399] = 3'b000;
        rom_memory[43400] = 3'b000;
        rom_memory[43401] = 3'b000;
        rom_memory[43402] = 3'b000;
        rom_memory[43403] = 3'b000;
        rom_memory[43404] = 3'b110;
        rom_memory[43405] = 3'b111;
        rom_memory[43406] = 3'b110;
        rom_memory[43407] = 3'b110;
        rom_memory[43408] = 3'b110;
        rom_memory[43409] = 3'b110;
        rom_memory[43410] = 3'b110;
        rom_memory[43411] = 3'b110;
        rom_memory[43412] = 3'b110;
        rom_memory[43413] = 3'b110;
        rom_memory[43414] = 3'b110;
        rom_memory[43415] = 3'b110;
        rom_memory[43416] = 3'b110;
        rom_memory[43417] = 3'b110;
        rom_memory[43418] = 3'b110;
        rom_memory[43419] = 3'b110;
        rom_memory[43420] = 3'b110;
        rom_memory[43421] = 3'b110;
        rom_memory[43422] = 3'b110;
        rom_memory[43423] = 3'b110;
        rom_memory[43424] = 3'b110;
        rom_memory[43425] = 3'b110;
        rom_memory[43426] = 3'b110;
        rom_memory[43427] = 3'b110;
        rom_memory[43428] = 3'b110;
        rom_memory[43429] = 3'b110;
        rom_memory[43430] = 3'b110;
        rom_memory[43431] = 3'b110;
        rom_memory[43432] = 3'b110;
        rom_memory[43433] = 3'b110;
        rom_memory[43434] = 3'b110;
        rom_memory[43435] = 3'b110;
        rom_memory[43436] = 3'b110;
        rom_memory[43437] = 3'b110;
        rom_memory[43438] = 3'b110;
        rom_memory[43439] = 3'b110;
        rom_memory[43440] = 3'b111;
        rom_memory[43441] = 3'b111;
        rom_memory[43442] = 3'b111;
        rom_memory[43443] = 3'b111;
        rom_memory[43444] = 3'b111;
        rom_memory[43445] = 3'b111;
        rom_memory[43446] = 3'b111;
        rom_memory[43447] = 3'b111;
        rom_memory[43448] = 3'b111;
        rom_memory[43449] = 3'b111;
        rom_memory[43450] = 3'b111;
        rom_memory[43451] = 3'b111;
        rom_memory[43452] = 3'b111;
        rom_memory[43453] = 3'b111;
        rom_memory[43454] = 3'b111;
        rom_memory[43455] = 3'b111;
        rom_memory[43456] = 3'b111;
        rom_memory[43457] = 3'b111;
        rom_memory[43458] = 3'b111;
        rom_memory[43459] = 3'b111;
        rom_memory[43460] = 3'b111;
        rom_memory[43461] = 3'b110;
        rom_memory[43462] = 3'b110;
        rom_memory[43463] = 3'b110;
        rom_memory[43464] = 3'b110;
        rom_memory[43465] = 3'b110;
        rom_memory[43466] = 3'b110;
        rom_memory[43467] = 3'b110;
        rom_memory[43468] = 3'b110;
        rom_memory[43469] = 3'b110;
        rom_memory[43470] = 3'b110;
        rom_memory[43471] = 3'b110;
        rom_memory[43472] = 3'b111;
        rom_memory[43473] = 3'b111;
        rom_memory[43474] = 3'b111;
        rom_memory[43475] = 3'b111;
        rom_memory[43476] = 3'b111;
        rom_memory[43477] = 3'b111;
        rom_memory[43478] = 3'b111;
        rom_memory[43479] = 3'b111;
        rom_memory[43480] = 3'b111;
        rom_memory[43481] = 3'b111;
        rom_memory[43482] = 3'b111;
        rom_memory[43483] = 3'b111;
        rom_memory[43484] = 3'b111;
        rom_memory[43485] = 3'b110;
        rom_memory[43486] = 3'b110;
        rom_memory[43487] = 3'b110;
        rom_memory[43488] = 3'b110;
        rom_memory[43489] = 3'b111;
        rom_memory[43490] = 3'b111;
        rom_memory[43491] = 3'b111;
        rom_memory[43492] = 3'b111;
        rom_memory[43493] = 3'b111;
        rom_memory[43494] = 3'b111;
        rom_memory[43495] = 3'b111;
        rom_memory[43496] = 3'b111;
        rom_memory[43497] = 3'b110;
        rom_memory[43498] = 3'b110;
        rom_memory[43499] = 3'b111;
        rom_memory[43500] = 3'b110;
        rom_memory[43501] = 3'b110;
        rom_memory[43502] = 3'b100;
        rom_memory[43503] = 3'b111;
        rom_memory[43504] = 3'b110;
        rom_memory[43505] = 3'b110;
        rom_memory[43506] = 3'b110;
        rom_memory[43507] = 3'b111;
        rom_memory[43508] = 3'b110;
        rom_memory[43509] = 3'b110;
        rom_memory[43510] = 3'b111;
        rom_memory[43511] = 3'b110;
        rom_memory[43512] = 3'b000;
        rom_memory[43513] = 3'b100;
        rom_memory[43514] = 3'b000;
        rom_memory[43515] = 3'b110;
        rom_memory[43516] = 3'b100;
        rom_memory[43517] = 3'b100;
        rom_memory[43518] = 3'b100;
        rom_memory[43519] = 3'b110;
        rom_memory[43520] = 3'b111;
        rom_memory[43521] = 3'b110;
        rom_memory[43522] = 3'b111;
        rom_memory[43523] = 3'b110;
        rom_memory[43524] = 3'b110;
        rom_memory[43525] = 3'b110;
        rom_memory[43526] = 3'b110;
        rom_memory[43527] = 3'b110;
        rom_memory[43528] = 3'b110;
        rom_memory[43529] = 3'b110;
        rom_memory[43530] = 3'b110;
        rom_memory[43531] = 3'b110;
        rom_memory[43532] = 3'b110;
        rom_memory[43533] = 3'b111;
        rom_memory[43534] = 3'b111;
        rom_memory[43535] = 3'b111;
        rom_memory[43536] = 3'b111;
        rom_memory[43537] = 3'b111;
        rom_memory[43538] = 3'b111;
        rom_memory[43539] = 3'b110;
        rom_memory[43540] = 3'b110;
        rom_memory[43541] = 3'b110;
        rom_memory[43542] = 3'b110;
        rom_memory[43543] = 3'b111;
        rom_memory[43544] = 3'b111;
        rom_memory[43545] = 3'b111;
        rom_memory[43546] = 3'b111;
        rom_memory[43547] = 3'b111;
        rom_memory[43548] = 3'b111;
        rom_memory[43549] = 3'b111;
        rom_memory[43550] = 3'b111;
        rom_memory[43551] = 3'b111;
        rom_memory[43552] = 3'b111;
        rom_memory[43553] = 3'b111;
        rom_memory[43554] = 3'b110;
        rom_memory[43555] = 3'b110;
        rom_memory[43556] = 3'b110;
        rom_memory[43557] = 3'b110;
        rom_memory[43558] = 3'b110;
        rom_memory[43559] = 3'b110;
        rom_memory[43560] = 3'b110;
        rom_memory[43561] = 3'b110;
        rom_memory[43562] = 3'b110;
        rom_memory[43563] = 3'b110;
        rom_memory[43564] = 3'b110;
        rom_memory[43565] = 3'b110;
        rom_memory[43566] = 3'b110;
        rom_memory[43567] = 3'b110;
        rom_memory[43568] = 3'b110;
        rom_memory[43569] = 3'b110;
        rom_memory[43570] = 3'b110;
        rom_memory[43571] = 3'b110;
        rom_memory[43572] = 3'b110;
        rom_memory[43573] = 3'b110;
        rom_memory[43574] = 3'b110;
        rom_memory[43575] = 3'b110;
        rom_memory[43576] = 3'b110;
        rom_memory[43577] = 3'b110;
        rom_memory[43578] = 3'b110;
        rom_memory[43579] = 3'b110;
        rom_memory[43580] = 3'b110;
        rom_memory[43581] = 3'b110;
        rom_memory[43582] = 3'b110;
        rom_memory[43583] = 3'b110;
        rom_memory[43584] = 3'b110;
        rom_memory[43585] = 3'b110;
        rom_memory[43586] = 3'b110;
        rom_memory[43587] = 3'b110;
        rom_memory[43588] = 3'b110;
        rom_memory[43589] = 3'b110;
        rom_memory[43590] = 3'b110;
        rom_memory[43591] = 3'b110;
        rom_memory[43592] = 3'b110;
        rom_memory[43593] = 3'b110;
        rom_memory[43594] = 3'b110;
        rom_memory[43595] = 3'b110;
        rom_memory[43596] = 3'b110;
        rom_memory[43597] = 3'b110;
        rom_memory[43598] = 3'b110;
        rom_memory[43599] = 3'b110;
        rom_memory[43600] = 3'b110;
        rom_memory[43601] = 3'b110;
        rom_memory[43602] = 3'b110;
        rom_memory[43603] = 3'b110;
        rom_memory[43604] = 3'b110;
        rom_memory[43605] = 3'b110;
        rom_memory[43606] = 3'b110;
        rom_memory[43607] = 3'b110;
        rom_memory[43608] = 3'b110;
        rom_memory[43609] = 3'b110;
        rom_memory[43610] = 3'b110;
        rom_memory[43611] = 3'b110;
        rom_memory[43612] = 3'b110;
        rom_memory[43613] = 3'b110;
        rom_memory[43614] = 3'b110;
        rom_memory[43615] = 3'b110;
        rom_memory[43616] = 3'b110;
        rom_memory[43617] = 3'b110;
        rom_memory[43618] = 3'b110;
        rom_memory[43619] = 3'b110;
        rom_memory[43620] = 3'b110;
        rom_memory[43621] = 3'b110;
        rom_memory[43622] = 3'b110;
        rom_memory[43623] = 3'b110;
        rom_memory[43624] = 3'b110;
        rom_memory[43625] = 3'b110;
        rom_memory[43626] = 3'b110;
        rom_memory[43627] = 3'b110;
        rom_memory[43628] = 3'b110;
        rom_memory[43629] = 3'b110;
        rom_memory[43630] = 3'b110;
        rom_memory[43631] = 3'b110;
        rom_memory[43632] = 3'b110;
        rom_memory[43633] = 3'b000;
        rom_memory[43634] = 3'b000;
        rom_memory[43635] = 3'b000;
        rom_memory[43636] = 3'b000;
        rom_memory[43637] = 3'b000;
        rom_memory[43638] = 3'b000;
        rom_memory[43639] = 3'b000;
        rom_memory[43640] = 3'b000;
        rom_memory[43641] = 3'b000;
        rom_memory[43642] = 3'b000;
        rom_memory[43643] = 3'b000;
        rom_memory[43644] = 3'b000;
        rom_memory[43645] = 3'b000;
        rom_memory[43646] = 3'b110;
        rom_memory[43647] = 3'b110;
        rom_memory[43648] = 3'b110;
        rom_memory[43649] = 3'b110;
        rom_memory[43650] = 3'b110;
        rom_memory[43651] = 3'b110;
        rom_memory[43652] = 3'b110;
        rom_memory[43653] = 3'b110;
        rom_memory[43654] = 3'b110;
        rom_memory[43655] = 3'b110;
        rom_memory[43656] = 3'b110;
        rom_memory[43657] = 3'b110;
        rom_memory[43658] = 3'b110;
        rom_memory[43659] = 3'b110;
        rom_memory[43660] = 3'b110;
        rom_memory[43661] = 3'b110;
        rom_memory[43662] = 3'b110;
        rom_memory[43663] = 3'b110;
        rom_memory[43664] = 3'b110;
        rom_memory[43665] = 3'b110;
        rom_memory[43666] = 3'b110;
        rom_memory[43667] = 3'b110;
        rom_memory[43668] = 3'b110;
        rom_memory[43669] = 3'b110;
        rom_memory[43670] = 3'b110;
        rom_memory[43671] = 3'b110;
        rom_memory[43672] = 3'b110;
        rom_memory[43673] = 3'b110;
        rom_memory[43674] = 3'b110;
        rom_memory[43675] = 3'b110;
        rom_memory[43676] = 3'b110;
        rom_memory[43677] = 3'b110;
        rom_memory[43678] = 3'b110;
        rom_memory[43679] = 3'b110;
        rom_memory[43680] = 3'b111;
        rom_memory[43681] = 3'b111;
        rom_memory[43682] = 3'b111;
        rom_memory[43683] = 3'b111;
        rom_memory[43684] = 3'b111;
        rom_memory[43685] = 3'b111;
        rom_memory[43686] = 3'b111;
        rom_memory[43687] = 3'b111;
        rom_memory[43688] = 3'b111;
        rom_memory[43689] = 3'b111;
        rom_memory[43690] = 3'b111;
        rom_memory[43691] = 3'b111;
        rom_memory[43692] = 3'b111;
        rom_memory[43693] = 3'b111;
        rom_memory[43694] = 3'b111;
        rom_memory[43695] = 3'b111;
        rom_memory[43696] = 3'b111;
        rom_memory[43697] = 3'b111;
        rom_memory[43698] = 3'b111;
        rom_memory[43699] = 3'b111;
        rom_memory[43700] = 3'b111;
        rom_memory[43701] = 3'b111;
        rom_memory[43702] = 3'b110;
        rom_memory[43703] = 3'b110;
        rom_memory[43704] = 3'b110;
        rom_memory[43705] = 3'b110;
        rom_memory[43706] = 3'b110;
        rom_memory[43707] = 3'b110;
        rom_memory[43708] = 3'b110;
        rom_memory[43709] = 3'b110;
        rom_memory[43710] = 3'b110;
        rom_memory[43711] = 3'b111;
        rom_memory[43712] = 3'b111;
        rom_memory[43713] = 3'b111;
        rom_memory[43714] = 3'b111;
        rom_memory[43715] = 3'b111;
        rom_memory[43716] = 3'b111;
        rom_memory[43717] = 3'b111;
        rom_memory[43718] = 3'b111;
        rom_memory[43719] = 3'b111;
        rom_memory[43720] = 3'b111;
        rom_memory[43721] = 3'b111;
        rom_memory[43722] = 3'b111;
        rom_memory[43723] = 3'b111;
        rom_memory[43724] = 3'b111;
        rom_memory[43725] = 3'b110;
        rom_memory[43726] = 3'b110;
        rom_memory[43727] = 3'b110;
        rom_memory[43728] = 3'b110;
        rom_memory[43729] = 3'b110;
        rom_memory[43730] = 3'b110;
        rom_memory[43731] = 3'b111;
        rom_memory[43732] = 3'b111;
        rom_memory[43733] = 3'b111;
        rom_memory[43734] = 3'b111;
        rom_memory[43735] = 3'b111;
        rom_memory[43736] = 3'b111;
        rom_memory[43737] = 3'b110;
        rom_memory[43738] = 3'b110;
        rom_memory[43739] = 3'b110;
        rom_memory[43740] = 3'b110;
        rom_memory[43741] = 3'b110;
        rom_memory[43742] = 3'b110;
        rom_memory[43743] = 3'b110;
        rom_memory[43744] = 3'b110;
        rom_memory[43745] = 3'b110;
        rom_memory[43746] = 3'b110;
        rom_memory[43747] = 3'b110;
        rom_memory[43748] = 3'b110;
        rom_memory[43749] = 3'b110;
        rom_memory[43750] = 3'b110;
        rom_memory[43751] = 3'b110;
        rom_memory[43752] = 3'b110;
        rom_memory[43753] = 3'b100;
        rom_memory[43754] = 3'b100;
        rom_memory[43755] = 3'b111;
        rom_memory[43756] = 3'b000;
        rom_memory[43757] = 3'b000;
        rom_memory[43758] = 3'b100;
        rom_memory[43759] = 3'b110;
        rom_memory[43760] = 3'b111;
        rom_memory[43761] = 3'b111;
        rom_memory[43762] = 3'b110;
        rom_memory[43763] = 3'b110;
        rom_memory[43764] = 3'b110;
        rom_memory[43765] = 3'b110;
        rom_memory[43766] = 3'b110;
        rom_memory[43767] = 3'b110;
        rom_memory[43768] = 3'b110;
        rom_memory[43769] = 3'b110;
        rom_memory[43770] = 3'b110;
        rom_memory[43771] = 3'b110;
        rom_memory[43772] = 3'b110;
        rom_memory[43773] = 3'b110;
        rom_memory[43774] = 3'b111;
        rom_memory[43775] = 3'b111;
        rom_memory[43776] = 3'b111;
        rom_memory[43777] = 3'b111;
        rom_memory[43778] = 3'b111;
        rom_memory[43779] = 3'b111;
        rom_memory[43780] = 3'b110;
        rom_memory[43781] = 3'b110;
        rom_memory[43782] = 3'b111;
        rom_memory[43783] = 3'b111;
        rom_memory[43784] = 3'b111;
        rom_memory[43785] = 3'b111;
        rom_memory[43786] = 3'b111;
        rom_memory[43787] = 3'b111;
        rom_memory[43788] = 3'b111;
        rom_memory[43789] = 3'b111;
        rom_memory[43790] = 3'b111;
        rom_memory[43791] = 3'b111;
        rom_memory[43792] = 3'b111;
        rom_memory[43793] = 3'b111;
        rom_memory[43794] = 3'b110;
        rom_memory[43795] = 3'b110;
        rom_memory[43796] = 3'b110;
        rom_memory[43797] = 3'b110;
        rom_memory[43798] = 3'b110;
        rom_memory[43799] = 3'b110;
        rom_memory[43800] = 3'b110;
        rom_memory[43801] = 3'b110;
        rom_memory[43802] = 3'b110;
        rom_memory[43803] = 3'b110;
        rom_memory[43804] = 3'b110;
        rom_memory[43805] = 3'b110;
        rom_memory[43806] = 3'b110;
        rom_memory[43807] = 3'b110;
        rom_memory[43808] = 3'b110;
        rom_memory[43809] = 3'b110;
        rom_memory[43810] = 3'b110;
        rom_memory[43811] = 3'b110;
        rom_memory[43812] = 3'b110;
        rom_memory[43813] = 3'b110;
        rom_memory[43814] = 3'b110;
        rom_memory[43815] = 3'b110;
        rom_memory[43816] = 3'b110;
        rom_memory[43817] = 3'b110;
        rom_memory[43818] = 3'b110;
        rom_memory[43819] = 3'b110;
        rom_memory[43820] = 3'b110;
        rom_memory[43821] = 3'b110;
        rom_memory[43822] = 3'b110;
        rom_memory[43823] = 3'b110;
        rom_memory[43824] = 3'b110;
        rom_memory[43825] = 3'b110;
        rom_memory[43826] = 3'b110;
        rom_memory[43827] = 3'b110;
        rom_memory[43828] = 3'b110;
        rom_memory[43829] = 3'b110;
        rom_memory[43830] = 3'b110;
        rom_memory[43831] = 3'b110;
        rom_memory[43832] = 3'b110;
        rom_memory[43833] = 3'b110;
        rom_memory[43834] = 3'b110;
        rom_memory[43835] = 3'b110;
        rom_memory[43836] = 3'b110;
        rom_memory[43837] = 3'b110;
        rom_memory[43838] = 3'b110;
        rom_memory[43839] = 3'b110;
        rom_memory[43840] = 3'b110;
        rom_memory[43841] = 3'b110;
        rom_memory[43842] = 3'b110;
        rom_memory[43843] = 3'b110;
        rom_memory[43844] = 3'b110;
        rom_memory[43845] = 3'b110;
        rom_memory[43846] = 3'b110;
        rom_memory[43847] = 3'b110;
        rom_memory[43848] = 3'b110;
        rom_memory[43849] = 3'b110;
        rom_memory[43850] = 3'b110;
        rom_memory[43851] = 3'b110;
        rom_memory[43852] = 3'b110;
        rom_memory[43853] = 3'b110;
        rom_memory[43854] = 3'b110;
        rom_memory[43855] = 3'b110;
        rom_memory[43856] = 3'b110;
        rom_memory[43857] = 3'b110;
        rom_memory[43858] = 3'b110;
        rom_memory[43859] = 3'b110;
        rom_memory[43860] = 3'b110;
        rom_memory[43861] = 3'b110;
        rom_memory[43862] = 3'b110;
        rom_memory[43863] = 3'b110;
        rom_memory[43864] = 3'b110;
        rom_memory[43865] = 3'b110;
        rom_memory[43866] = 3'b110;
        rom_memory[43867] = 3'b110;
        rom_memory[43868] = 3'b110;
        rom_memory[43869] = 3'b110;
        rom_memory[43870] = 3'b110;
        rom_memory[43871] = 3'b110;
        rom_memory[43872] = 3'b110;
        rom_memory[43873] = 3'b110;
        rom_memory[43874] = 3'b100;
        rom_memory[43875] = 3'b000;
        rom_memory[43876] = 3'b000;
        rom_memory[43877] = 3'b000;
        rom_memory[43878] = 3'b000;
        rom_memory[43879] = 3'b000;
        rom_memory[43880] = 3'b000;
        rom_memory[43881] = 3'b000;
        rom_memory[43882] = 3'b000;
        rom_memory[43883] = 3'b000;
        rom_memory[43884] = 3'b000;
        rom_memory[43885] = 3'b000;
        rom_memory[43886] = 3'b000;
        rom_memory[43887] = 3'b000;
        rom_memory[43888] = 3'b110;
        rom_memory[43889] = 3'b110;
        rom_memory[43890] = 3'b110;
        rom_memory[43891] = 3'b110;
        rom_memory[43892] = 3'b110;
        rom_memory[43893] = 3'b110;
        rom_memory[43894] = 3'b110;
        rom_memory[43895] = 3'b110;
        rom_memory[43896] = 3'b110;
        rom_memory[43897] = 3'b110;
        rom_memory[43898] = 3'b110;
        rom_memory[43899] = 3'b110;
        rom_memory[43900] = 3'b110;
        rom_memory[43901] = 3'b110;
        rom_memory[43902] = 3'b110;
        rom_memory[43903] = 3'b110;
        rom_memory[43904] = 3'b110;
        rom_memory[43905] = 3'b110;
        rom_memory[43906] = 3'b110;
        rom_memory[43907] = 3'b110;
        rom_memory[43908] = 3'b110;
        rom_memory[43909] = 3'b110;
        rom_memory[43910] = 3'b110;
        rom_memory[43911] = 3'b110;
        rom_memory[43912] = 3'b110;
        rom_memory[43913] = 3'b110;
        rom_memory[43914] = 3'b110;
        rom_memory[43915] = 3'b110;
        rom_memory[43916] = 3'b110;
        rom_memory[43917] = 3'b110;
        rom_memory[43918] = 3'b110;
        rom_memory[43919] = 3'b110;
        rom_memory[43920] = 3'b111;
        rom_memory[43921] = 3'b111;
        rom_memory[43922] = 3'b111;
        rom_memory[43923] = 3'b111;
        rom_memory[43924] = 3'b111;
        rom_memory[43925] = 3'b111;
        rom_memory[43926] = 3'b111;
        rom_memory[43927] = 3'b111;
        rom_memory[43928] = 3'b111;
        rom_memory[43929] = 3'b111;
        rom_memory[43930] = 3'b111;
        rom_memory[43931] = 3'b111;
        rom_memory[43932] = 3'b111;
        rom_memory[43933] = 3'b111;
        rom_memory[43934] = 3'b111;
        rom_memory[43935] = 3'b111;
        rom_memory[43936] = 3'b111;
        rom_memory[43937] = 3'b111;
        rom_memory[43938] = 3'b111;
        rom_memory[43939] = 3'b111;
        rom_memory[43940] = 3'b111;
        rom_memory[43941] = 3'b110;
        rom_memory[43942] = 3'b110;
        rom_memory[43943] = 3'b110;
        rom_memory[43944] = 3'b110;
        rom_memory[43945] = 3'b110;
        rom_memory[43946] = 3'b110;
        rom_memory[43947] = 3'b110;
        rom_memory[43948] = 3'b110;
        rom_memory[43949] = 3'b110;
        rom_memory[43950] = 3'b110;
        rom_memory[43951] = 3'b111;
        rom_memory[43952] = 3'b111;
        rom_memory[43953] = 3'b111;
        rom_memory[43954] = 3'b111;
        rom_memory[43955] = 3'b111;
        rom_memory[43956] = 3'b111;
        rom_memory[43957] = 3'b111;
        rom_memory[43958] = 3'b111;
        rom_memory[43959] = 3'b111;
        rom_memory[43960] = 3'b111;
        rom_memory[43961] = 3'b111;
        rom_memory[43962] = 3'b111;
        rom_memory[43963] = 3'b111;
        rom_memory[43964] = 3'b111;
        rom_memory[43965] = 3'b111;
        rom_memory[43966] = 3'b110;
        rom_memory[43967] = 3'b110;
        rom_memory[43968] = 3'b110;
        rom_memory[43969] = 3'b110;
        rom_memory[43970] = 3'b110;
        rom_memory[43971] = 3'b110;
        rom_memory[43972] = 3'b110;
        rom_memory[43973] = 3'b111;
        rom_memory[43974] = 3'b111;
        rom_memory[43975] = 3'b110;
        rom_memory[43976] = 3'b110;
        rom_memory[43977] = 3'b110;
        rom_memory[43978] = 3'b110;
        rom_memory[43979] = 3'b110;
        rom_memory[43980] = 3'b100;
        rom_memory[43981] = 3'b110;
        rom_memory[43982] = 3'b110;
        rom_memory[43983] = 3'b110;
        rom_memory[43984] = 3'b110;
        rom_memory[43985] = 3'b110;
        rom_memory[43986] = 3'b111;
        rom_memory[43987] = 3'b111;
        rom_memory[43988] = 3'b110;
        rom_memory[43989] = 3'b110;
        rom_memory[43990] = 3'b110;
        rom_memory[43991] = 3'b111;
        rom_memory[43992] = 3'b111;
        rom_memory[43993] = 3'b000;
        rom_memory[43994] = 3'b100;
        rom_memory[43995] = 3'b000;
        rom_memory[43996] = 3'b000;
        rom_memory[43997] = 3'b000;
        rom_memory[43998] = 3'b000;
        rom_memory[43999] = 3'b111;
        rom_memory[44000] = 3'b111;
        rom_memory[44001] = 3'b110;
        rom_memory[44002] = 3'b110;
        rom_memory[44003] = 3'b110;
        rom_memory[44004] = 3'b110;
        rom_memory[44005] = 3'b110;
        rom_memory[44006] = 3'b110;
        rom_memory[44007] = 3'b110;
        rom_memory[44008] = 3'b110;
        rom_memory[44009] = 3'b110;
        rom_memory[44010] = 3'b110;
        rom_memory[44011] = 3'b110;
        rom_memory[44012] = 3'b110;
        rom_memory[44013] = 3'b110;
        rom_memory[44014] = 3'b111;
        rom_memory[44015] = 3'b111;
        rom_memory[44016] = 3'b111;
        rom_memory[44017] = 3'b111;
        rom_memory[44018] = 3'b111;
        rom_memory[44019] = 3'b111;
        rom_memory[44020] = 3'b111;
        rom_memory[44021] = 3'b111;
        rom_memory[44022] = 3'b111;
        rom_memory[44023] = 3'b111;
        rom_memory[44024] = 3'b111;
        rom_memory[44025] = 3'b111;
        rom_memory[44026] = 3'b111;
        rom_memory[44027] = 3'b111;
        rom_memory[44028] = 3'b111;
        rom_memory[44029] = 3'b111;
        rom_memory[44030] = 3'b111;
        rom_memory[44031] = 3'b111;
        rom_memory[44032] = 3'b111;
        rom_memory[44033] = 3'b111;
        rom_memory[44034] = 3'b110;
        rom_memory[44035] = 3'b110;
        rom_memory[44036] = 3'b110;
        rom_memory[44037] = 3'b110;
        rom_memory[44038] = 3'b110;
        rom_memory[44039] = 3'b110;
        rom_memory[44040] = 3'b110;
        rom_memory[44041] = 3'b110;
        rom_memory[44042] = 3'b110;
        rom_memory[44043] = 3'b110;
        rom_memory[44044] = 3'b110;
        rom_memory[44045] = 3'b110;
        rom_memory[44046] = 3'b110;
        rom_memory[44047] = 3'b110;
        rom_memory[44048] = 3'b110;
        rom_memory[44049] = 3'b110;
        rom_memory[44050] = 3'b110;
        rom_memory[44051] = 3'b110;
        rom_memory[44052] = 3'b110;
        rom_memory[44053] = 3'b110;
        rom_memory[44054] = 3'b110;
        rom_memory[44055] = 3'b110;
        rom_memory[44056] = 3'b110;
        rom_memory[44057] = 3'b110;
        rom_memory[44058] = 3'b110;
        rom_memory[44059] = 3'b110;
        rom_memory[44060] = 3'b110;
        rom_memory[44061] = 3'b110;
        rom_memory[44062] = 3'b110;
        rom_memory[44063] = 3'b110;
        rom_memory[44064] = 3'b110;
        rom_memory[44065] = 3'b110;
        rom_memory[44066] = 3'b110;
        rom_memory[44067] = 3'b110;
        rom_memory[44068] = 3'b110;
        rom_memory[44069] = 3'b110;
        rom_memory[44070] = 3'b110;
        rom_memory[44071] = 3'b110;
        rom_memory[44072] = 3'b110;
        rom_memory[44073] = 3'b110;
        rom_memory[44074] = 3'b110;
        rom_memory[44075] = 3'b110;
        rom_memory[44076] = 3'b110;
        rom_memory[44077] = 3'b110;
        rom_memory[44078] = 3'b110;
        rom_memory[44079] = 3'b110;
        rom_memory[44080] = 3'b110;
        rom_memory[44081] = 3'b110;
        rom_memory[44082] = 3'b110;
        rom_memory[44083] = 3'b110;
        rom_memory[44084] = 3'b110;
        rom_memory[44085] = 3'b110;
        rom_memory[44086] = 3'b110;
        rom_memory[44087] = 3'b110;
        rom_memory[44088] = 3'b110;
        rom_memory[44089] = 3'b110;
        rom_memory[44090] = 3'b110;
        rom_memory[44091] = 3'b110;
        rom_memory[44092] = 3'b110;
        rom_memory[44093] = 3'b110;
        rom_memory[44094] = 3'b110;
        rom_memory[44095] = 3'b110;
        rom_memory[44096] = 3'b110;
        rom_memory[44097] = 3'b110;
        rom_memory[44098] = 3'b110;
        rom_memory[44099] = 3'b110;
        rom_memory[44100] = 3'b110;
        rom_memory[44101] = 3'b110;
        rom_memory[44102] = 3'b110;
        rom_memory[44103] = 3'b110;
        rom_memory[44104] = 3'b110;
        rom_memory[44105] = 3'b110;
        rom_memory[44106] = 3'b110;
        rom_memory[44107] = 3'b110;
        rom_memory[44108] = 3'b110;
        rom_memory[44109] = 3'b110;
        rom_memory[44110] = 3'b110;
        rom_memory[44111] = 3'b110;
        rom_memory[44112] = 3'b110;
        rom_memory[44113] = 3'b110;
        rom_memory[44114] = 3'b110;
        rom_memory[44115] = 3'b110;
        rom_memory[44116] = 3'b100;
        rom_memory[44117] = 3'b000;
        rom_memory[44118] = 3'b000;
        rom_memory[44119] = 3'b000;
        rom_memory[44120] = 3'b000;
        rom_memory[44121] = 3'b000;
        rom_memory[44122] = 3'b000;
        rom_memory[44123] = 3'b000;
        rom_memory[44124] = 3'b100;
        rom_memory[44125] = 3'b100;
        rom_memory[44126] = 3'b000;
        rom_memory[44127] = 3'b000;
        rom_memory[44128] = 3'b000;
        rom_memory[44129] = 3'b000;
        rom_memory[44130] = 3'b110;
        rom_memory[44131] = 3'b110;
        rom_memory[44132] = 3'b110;
        rom_memory[44133] = 3'b110;
        rom_memory[44134] = 3'b110;
        rom_memory[44135] = 3'b110;
        rom_memory[44136] = 3'b110;
        rom_memory[44137] = 3'b110;
        rom_memory[44138] = 3'b110;
        rom_memory[44139] = 3'b110;
        rom_memory[44140] = 3'b110;
        rom_memory[44141] = 3'b110;
        rom_memory[44142] = 3'b110;
        rom_memory[44143] = 3'b110;
        rom_memory[44144] = 3'b110;
        rom_memory[44145] = 3'b110;
        rom_memory[44146] = 3'b110;
        rom_memory[44147] = 3'b110;
        rom_memory[44148] = 3'b110;
        rom_memory[44149] = 3'b110;
        rom_memory[44150] = 3'b110;
        rom_memory[44151] = 3'b110;
        rom_memory[44152] = 3'b110;
        rom_memory[44153] = 3'b110;
        rom_memory[44154] = 3'b110;
        rom_memory[44155] = 3'b110;
        rom_memory[44156] = 3'b110;
        rom_memory[44157] = 3'b110;
        rom_memory[44158] = 3'b110;
        rom_memory[44159] = 3'b110;
        rom_memory[44160] = 3'b111;
        rom_memory[44161] = 3'b111;
        rom_memory[44162] = 3'b111;
        rom_memory[44163] = 3'b111;
        rom_memory[44164] = 3'b111;
        rom_memory[44165] = 3'b111;
        rom_memory[44166] = 3'b111;
        rom_memory[44167] = 3'b111;
        rom_memory[44168] = 3'b111;
        rom_memory[44169] = 3'b111;
        rom_memory[44170] = 3'b111;
        rom_memory[44171] = 3'b111;
        rom_memory[44172] = 3'b111;
        rom_memory[44173] = 3'b111;
        rom_memory[44174] = 3'b111;
        rom_memory[44175] = 3'b111;
        rom_memory[44176] = 3'b111;
        rom_memory[44177] = 3'b111;
        rom_memory[44178] = 3'b111;
        rom_memory[44179] = 3'b111;
        rom_memory[44180] = 3'b111;
        rom_memory[44181] = 3'b110;
        rom_memory[44182] = 3'b110;
        rom_memory[44183] = 3'b110;
        rom_memory[44184] = 3'b110;
        rom_memory[44185] = 3'b110;
        rom_memory[44186] = 3'b110;
        rom_memory[44187] = 3'b110;
        rom_memory[44188] = 3'b110;
        rom_memory[44189] = 3'b110;
        rom_memory[44190] = 3'b110;
        rom_memory[44191] = 3'b111;
        rom_memory[44192] = 3'b111;
        rom_memory[44193] = 3'b111;
        rom_memory[44194] = 3'b111;
        rom_memory[44195] = 3'b111;
        rom_memory[44196] = 3'b111;
        rom_memory[44197] = 3'b111;
        rom_memory[44198] = 3'b111;
        rom_memory[44199] = 3'b111;
        rom_memory[44200] = 3'b111;
        rom_memory[44201] = 3'b111;
        rom_memory[44202] = 3'b111;
        rom_memory[44203] = 3'b111;
        rom_memory[44204] = 3'b111;
        rom_memory[44205] = 3'b111;
        rom_memory[44206] = 3'b111;
        rom_memory[44207] = 3'b111;
        rom_memory[44208] = 3'b110;
        rom_memory[44209] = 3'b110;
        rom_memory[44210] = 3'b110;
        rom_memory[44211] = 3'b110;
        rom_memory[44212] = 3'b110;
        rom_memory[44213] = 3'b110;
        rom_memory[44214] = 3'b110;
        rom_memory[44215] = 3'b110;
        rom_memory[44216] = 3'b110;
        rom_memory[44217] = 3'b110;
        rom_memory[44218] = 3'b100;
        rom_memory[44219] = 3'b110;
        rom_memory[44220] = 3'b100;
        rom_memory[44221] = 3'b100;
        rom_memory[44222] = 3'b110;
        rom_memory[44223] = 3'b100;
        rom_memory[44224] = 3'b110;
        rom_memory[44225] = 3'b110;
        rom_memory[44226] = 3'b111;
        rom_memory[44227] = 3'b111;
        rom_memory[44228] = 3'b110;
        rom_memory[44229] = 3'b110;
        rom_memory[44230] = 3'b110;
        rom_memory[44231] = 3'b110;
        rom_memory[44232] = 3'b111;
        rom_memory[44233] = 3'b100;
        rom_memory[44234] = 3'b000;
        rom_memory[44235] = 3'b000;
        rom_memory[44236] = 3'b000;
        rom_memory[44237] = 3'b000;
        rom_memory[44238] = 3'b000;
        rom_memory[44239] = 3'b100;
        rom_memory[44240] = 3'b111;
        rom_memory[44241] = 3'b110;
        rom_memory[44242] = 3'b110;
        rom_memory[44243] = 3'b110;
        rom_memory[44244] = 3'b110;
        rom_memory[44245] = 3'b111;
        rom_memory[44246] = 3'b111;
        rom_memory[44247] = 3'b110;
        rom_memory[44248] = 3'b110;
        rom_memory[44249] = 3'b110;
        rom_memory[44250] = 3'b110;
        rom_memory[44251] = 3'b110;
        rom_memory[44252] = 3'b110;
        rom_memory[44253] = 3'b110;
        rom_memory[44254] = 3'b110;
        rom_memory[44255] = 3'b110;
        rom_memory[44256] = 3'b110;
        rom_memory[44257] = 3'b111;
        rom_memory[44258] = 3'b111;
        rom_memory[44259] = 3'b111;
        rom_memory[44260] = 3'b111;
        rom_memory[44261] = 3'b111;
        rom_memory[44262] = 3'b111;
        rom_memory[44263] = 3'b111;
        rom_memory[44264] = 3'b111;
        rom_memory[44265] = 3'b111;
        rom_memory[44266] = 3'b111;
        rom_memory[44267] = 3'b111;
        rom_memory[44268] = 3'b111;
        rom_memory[44269] = 3'b111;
        rom_memory[44270] = 3'b111;
        rom_memory[44271] = 3'b111;
        rom_memory[44272] = 3'b111;
        rom_memory[44273] = 3'b111;
        rom_memory[44274] = 3'b111;
        rom_memory[44275] = 3'b110;
        rom_memory[44276] = 3'b110;
        rom_memory[44277] = 3'b110;
        rom_memory[44278] = 3'b110;
        rom_memory[44279] = 3'b110;
        rom_memory[44280] = 3'b110;
        rom_memory[44281] = 3'b110;
        rom_memory[44282] = 3'b110;
        rom_memory[44283] = 3'b110;
        rom_memory[44284] = 3'b110;
        rom_memory[44285] = 3'b110;
        rom_memory[44286] = 3'b110;
        rom_memory[44287] = 3'b110;
        rom_memory[44288] = 3'b110;
        rom_memory[44289] = 3'b110;
        rom_memory[44290] = 3'b110;
        rom_memory[44291] = 3'b110;
        rom_memory[44292] = 3'b110;
        rom_memory[44293] = 3'b110;
        rom_memory[44294] = 3'b110;
        rom_memory[44295] = 3'b110;
        rom_memory[44296] = 3'b110;
        rom_memory[44297] = 3'b110;
        rom_memory[44298] = 3'b110;
        rom_memory[44299] = 3'b110;
        rom_memory[44300] = 3'b110;
        rom_memory[44301] = 3'b110;
        rom_memory[44302] = 3'b110;
        rom_memory[44303] = 3'b110;
        rom_memory[44304] = 3'b110;
        rom_memory[44305] = 3'b110;
        rom_memory[44306] = 3'b110;
        rom_memory[44307] = 3'b110;
        rom_memory[44308] = 3'b110;
        rom_memory[44309] = 3'b110;
        rom_memory[44310] = 3'b110;
        rom_memory[44311] = 3'b110;
        rom_memory[44312] = 3'b110;
        rom_memory[44313] = 3'b110;
        rom_memory[44314] = 3'b110;
        rom_memory[44315] = 3'b110;
        rom_memory[44316] = 3'b110;
        rom_memory[44317] = 3'b110;
        rom_memory[44318] = 3'b110;
        rom_memory[44319] = 3'b110;
        rom_memory[44320] = 3'b110;
        rom_memory[44321] = 3'b110;
        rom_memory[44322] = 3'b110;
        rom_memory[44323] = 3'b110;
        rom_memory[44324] = 3'b110;
        rom_memory[44325] = 3'b110;
        rom_memory[44326] = 3'b110;
        rom_memory[44327] = 3'b110;
        rom_memory[44328] = 3'b110;
        rom_memory[44329] = 3'b110;
        rom_memory[44330] = 3'b110;
        rom_memory[44331] = 3'b110;
        rom_memory[44332] = 3'b110;
        rom_memory[44333] = 3'b110;
        rom_memory[44334] = 3'b110;
        rom_memory[44335] = 3'b110;
        rom_memory[44336] = 3'b110;
        rom_memory[44337] = 3'b110;
        rom_memory[44338] = 3'b110;
        rom_memory[44339] = 3'b110;
        rom_memory[44340] = 3'b110;
        rom_memory[44341] = 3'b110;
        rom_memory[44342] = 3'b110;
        rom_memory[44343] = 3'b110;
        rom_memory[44344] = 3'b110;
        rom_memory[44345] = 3'b110;
        rom_memory[44346] = 3'b110;
        rom_memory[44347] = 3'b110;
        rom_memory[44348] = 3'b110;
        rom_memory[44349] = 3'b110;
        rom_memory[44350] = 3'b110;
        rom_memory[44351] = 3'b110;
        rom_memory[44352] = 3'b110;
        rom_memory[44353] = 3'b110;
        rom_memory[44354] = 3'b110;
        rom_memory[44355] = 3'b110;
        rom_memory[44356] = 3'b110;
        rom_memory[44357] = 3'b110;
        rom_memory[44358] = 3'b000;
        rom_memory[44359] = 3'b000;
        rom_memory[44360] = 3'b000;
        rom_memory[44361] = 3'b000;
        rom_memory[44362] = 3'b000;
        rom_memory[44363] = 3'b000;
        rom_memory[44364] = 3'b000;
        rom_memory[44365] = 3'b000;
        rom_memory[44366] = 3'b110;
        rom_memory[44367] = 3'b110;
        rom_memory[44368] = 3'b000;
        rom_memory[44369] = 3'b000;
        rom_memory[44370] = 3'b000;
        rom_memory[44371] = 3'b000;
        rom_memory[44372] = 3'b110;
        rom_memory[44373] = 3'b110;
        rom_memory[44374] = 3'b110;
        rom_memory[44375] = 3'b110;
        rom_memory[44376] = 3'b110;
        rom_memory[44377] = 3'b110;
        rom_memory[44378] = 3'b110;
        rom_memory[44379] = 3'b110;
        rom_memory[44380] = 3'b110;
        rom_memory[44381] = 3'b110;
        rom_memory[44382] = 3'b110;
        rom_memory[44383] = 3'b110;
        rom_memory[44384] = 3'b110;
        rom_memory[44385] = 3'b110;
        rom_memory[44386] = 3'b110;
        rom_memory[44387] = 3'b110;
        rom_memory[44388] = 3'b110;
        rom_memory[44389] = 3'b110;
        rom_memory[44390] = 3'b110;
        rom_memory[44391] = 3'b110;
        rom_memory[44392] = 3'b110;
        rom_memory[44393] = 3'b110;
        rom_memory[44394] = 3'b110;
        rom_memory[44395] = 3'b110;
        rom_memory[44396] = 3'b110;
        rom_memory[44397] = 3'b110;
        rom_memory[44398] = 3'b110;
        rom_memory[44399] = 3'b110;
        rom_memory[44400] = 3'b111;
        rom_memory[44401] = 3'b111;
        rom_memory[44402] = 3'b111;
        rom_memory[44403] = 3'b111;
        rom_memory[44404] = 3'b111;
        rom_memory[44405] = 3'b111;
        rom_memory[44406] = 3'b111;
        rom_memory[44407] = 3'b111;
        rom_memory[44408] = 3'b111;
        rom_memory[44409] = 3'b111;
        rom_memory[44410] = 3'b111;
        rom_memory[44411] = 3'b111;
        rom_memory[44412] = 3'b111;
        rom_memory[44413] = 3'b111;
        rom_memory[44414] = 3'b111;
        rom_memory[44415] = 3'b111;
        rom_memory[44416] = 3'b111;
        rom_memory[44417] = 3'b111;
        rom_memory[44418] = 3'b111;
        rom_memory[44419] = 3'b111;
        rom_memory[44420] = 3'b111;
        rom_memory[44421] = 3'b111;
        rom_memory[44422] = 3'b110;
        rom_memory[44423] = 3'b110;
        rom_memory[44424] = 3'b110;
        rom_memory[44425] = 3'b110;
        rom_memory[44426] = 3'b110;
        rom_memory[44427] = 3'b110;
        rom_memory[44428] = 3'b110;
        rom_memory[44429] = 3'b110;
        rom_memory[44430] = 3'b110;
        rom_memory[44431] = 3'b111;
        rom_memory[44432] = 3'b111;
        rom_memory[44433] = 3'b111;
        rom_memory[44434] = 3'b111;
        rom_memory[44435] = 3'b111;
        rom_memory[44436] = 3'b111;
        rom_memory[44437] = 3'b111;
        rom_memory[44438] = 3'b111;
        rom_memory[44439] = 3'b111;
        rom_memory[44440] = 3'b111;
        rom_memory[44441] = 3'b111;
        rom_memory[44442] = 3'b111;
        rom_memory[44443] = 3'b111;
        rom_memory[44444] = 3'b111;
        rom_memory[44445] = 3'b111;
        rom_memory[44446] = 3'b111;
        rom_memory[44447] = 3'b111;
        rom_memory[44448] = 3'b111;
        rom_memory[44449] = 3'b111;
        rom_memory[44450] = 3'b111;
        rom_memory[44451] = 3'b111;
        rom_memory[44452] = 3'b111;
        rom_memory[44453] = 3'b111;
        rom_memory[44454] = 3'b110;
        rom_memory[44455] = 3'b110;
        rom_memory[44456] = 3'b110;
        rom_memory[44457] = 3'b100;
        rom_memory[44458] = 3'b100;
        rom_memory[44459] = 3'b100;
        rom_memory[44460] = 3'b110;
        rom_memory[44461] = 3'b100;
        rom_memory[44462] = 3'b110;
        rom_memory[44463] = 3'b100;
        rom_memory[44464] = 3'b110;
        rom_memory[44465] = 3'b110;
        rom_memory[44466] = 3'b111;
        rom_memory[44467] = 3'b111;
        rom_memory[44468] = 3'b111;
        rom_memory[44469] = 3'b110;
        rom_memory[44470] = 3'b110;
        rom_memory[44471] = 3'b111;
        rom_memory[44472] = 3'b111;
        rom_memory[44473] = 3'b111;
        rom_memory[44474] = 3'b000;
        rom_memory[44475] = 3'b000;
        rom_memory[44476] = 3'b000;
        rom_memory[44477] = 3'b000;
        rom_memory[44478] = 3'b100;
        rom_memory[44479] = 3'b110;
        rom_memory[44480] = 3'b110;
        rom_memory[44481] = 3'b110;
        rom_memory[44482] = 3'b110;
        rom_memory[44483] = 3'b110;
        rom_memory[44484] = 3'b111;
        rom_memory[44485] = 3'b111;
        rom_memory[44486] = 3'b111;
        rom_memory[44487] = 3'b110;
        rom_memory[44488] = 3'b110;
        rom_memory[44489] = 3'b110;
        rom_memory[44490] = 3'b110;
        rom_memory[44491] = 3'b110;
        rom_memory[44492] = 3'b110;
        rom_memory[44493] = 3'b110;
        rom_memory[44494] = 3'b110;
        rom_memory[44495] = 3'b110;
        rom_memory[44496] = 3'b110;
        rom_memory[44497] = 3'b110;
        rom_memory[44498] = 3'b110;
        rom_memory[44499] = 3'b111;
        rom_memory[44500] = 3'b111;
        rom_memory[44501] = 3'b111;
        rom_memory[44502] = 3'b111;
        rom_memory[44503] = 3'b111;
        rom_memory[44504] = 3'b111;
        rom_memory[44505] = 3'b111;
        rom_memory[44506] = 3'b111;
        rom_memory[44507] = 3'b111;
        rom_memory[44508] = 3'b111;
        rom_memory[44509] = 3'b111;
        rom_memory[44510] = 3'b111;
        rom_memory[44511] = 3'b111;
        rom_memory[44512] = 3'b111;
        rom_memory[44513] = 3'b111;
        rom_memory[44514] = 3'b111;
        rom_memory[44515] = 3'b110;
        rom_memory[44516] = 3'b110;
        rom_memory[44517] = 3'b110;
        rom_memory[44518] = 3'b110;
        rom_memory[44519] = 3'b110;
        rom_memory[44520] = 3'b110;
        rom_memory[44521] = 3'b110;
        rom_memory[44522] = 3'b110;
        rom_memory[44523] = 3'b110;
        rom_memory[44524] = 3'b110;
        rom_memory[44525] = 3'b110;
        rom_memory[44526] = 3'b110;
        rom_memory[44527] = 3'b110;
        rom_memory[44528] = 3'b110;
        rom_memory[44529] = 3'b110;
        rom_memory[44530] = 3'b110;
        rom_memory[44531] = 3'b110;
        rom_memory[44532] = 3'b110;
        rom_memory[44533] = 3'b110;
        rom_memory[44534] = 3'b110;
        rom_memory[44535] = 3'b110;
        rom_memory[44536] = 3'b110;
        rom_memory[44537] = 3'b110;
        rom_memory[44538] = 3'b110;
        rom_memory[44539] = 3'b110;
        rom_memory[44540] = 3'b110;
        rom_memory[44541] = 3'b110;
        rom_memory[44542] = 3'b110;
        rom_memory[44543] = 3'b110;
        rom_memory[44544] = 3'b110;
        rom_memory[44545] = 3'b110;
        rom_memory[44546] = 3'b110;
        rom_memory[44547] = 3'b110;
        rom_memory[44548] = 3'b110;
        rom_memory[44549] = 3'b110;
        rom_memory[44550] = 3'b110;
        rom_memory[44551] = 3'b110;
        rom_memory[44552] = 3'b110;
        rom_memory[44553] = 3'b110;
        rom_memory[44554] = 3'b110;
        rom_memory[44555] = 3'b110;
        rom_memory[44556] = 3'b110;
        rom_memory[44557] = 3'b110;
        rom_memory[44558] = 3'b110;
        rom_memory[44559] = 3'b110;
        rom_memory[44560] = 3'b110;
        rom_memory[44561] = 3'b110;
        rom_memory[44562] = 3'b110;
        rom_memory[44563] = 3'b110;
        rom_memory[44564] = 3'b110;
        rom_memory[44565] = 3'b110;
        rom_memory[44566] = 3'b110;
        rom_memory[44567] = 3'b110;
        rom_memory[44568] = 3'b110;
        rom_memory[44569] = 3'b110;
        rom_memory[44570] = 3'b110;
        rom_memory[44571] = 3'b110;
        rom_memory[44572] = 3'b110;
        rom_memory[44573] = 3'b110;
        rom_memory[44574] = 3'b110;
        rom_memory[44575] = 3'b110;
        rom_memory[44576] = 3'b110;
        rom_memory[44577] = 3'b110;
        rom_memory[44578] = 3'b110;
        rom_memory[44579] = 3'b110;
        rom_memory[44580] = 3'b110;
        rom_memory[44581] = 3'b110;
        rom_memory[44582] = 3'b110;
        rom_memory[44583] = 3'b110;
        rom_memory[44584] = 3'b110;
        rom_memory[44585] = 3'b110;
        rom_memory[44586] = 3'b110;
        rom_memory[44587] = 3'b110;
        rom_memory[44588] = 3'b110;
        rom_memory[44589] = 3'b110;
        rom_memory[44590] = 3'b110;
        rom_memory[44591] = 3'b110;
        rom_memory[44592] = 3'b110;
        rom_memory[44593] = 3'b110;
        rom_memory[44594] = 3'b110;
        rom_memory[44595] = 3'b110;
        rom_memory[44596] = 3'b110;
        rom_memory[44597] = 3'b110;
        rom_memory[44598] = 3'b110;
        rom_memory[44599] = 3'b100;
        rom_memory[44600] = 3'b000;
        rom_memory[44601] = 3'b000;
        rom_memory[44602] = 3'b000;
        rom_memory[44603] = 3'b000;
        rom_memory[44604] = 3'b000;
        rom_memory[44605] = 3'b000;
        rom_memory[44606] = 3'b000;
        rom_memory[44607] = 3'b110;
        rom_memory[44608] = 3'b110;
        rom_memory[44609] = 3'b110;
        rom_memory[44610] = 3'b100;
        rom_memory[44611] = 3'b000;
        rom_memory[44612] = 3'b000;
        rom_memory[44613] = 3'b000;
        rom_memory[44614] = 3'b110;
        rom_memory[44615] = 3'b110;
        rom_memory[44616] = 3'b110;
        rom_memory[44617] = 3'b110;
        rom_memory[44618] = 3'b110;
        rom_memory[44619] = 3'b110;
        rom_memory[44620] = 3'b110;
        rom_memory[44621] = 3'b110;
        rom_memory[44622] = 3'b110;
        rom_memory[44623] = 3'b110;
        rom_memory[44624] = 3'b110;
        rom_memory[44625] = 3'b110;
        rom_memory[44626] = 3'b110;
        rom_memory[44627] = 3'b110;
        rom_memory[44628] = 3'b110;
        rom_memory[44629] = 3'b110;
        rom_memory[44630] = 3'b110;
        rom_memory[44631] = 3'b110;
        rom_memory[44632] = 3'b110;
        rom_memory[44633] = 3'b110;
        rom_memory[44634] = 3'b110;
        rom_memory[44635] = 3'b110;
        rom_memory[44636] = 3'b110;
        rom_memory[44637] = 3'b110;
        rom_memory[44638] = 3'b110;
        rom_memory[44639] = 3'b110;
        rom_memory[44640] = 3'b111;
        rom_memory[44641] = 3'b111;
        rom_memory[44642] = 3'b111;
        rom_memory[44643] = 3'b111;
        rom_memory[44644] = 3'b111;
        rom_memory[44645] = 3'b111;
        rom_memory[44646] = 3'b111;
        rom_memory[44647] = 3'b111;
        rom_memory[44648] = 3'b111;
        rom_memory[44649] = 3'b111;
        rom_memory[44650] = 3'b111;
        rom_memory[44651] = 3'b111;
        rom_memory[44652] = 3'b111;
        rom_memory[44653] = 3'b111;
        rom_memory[44654] = 3'b111;
        rom_memory[44655] = 3'b111;
        rom_memory[44656] = 3'b111;
        rom_memory[44657] = 3'b111;
        rom_memory[44658] = 3'b111;
        rom_memory[44659] = 3'b111;
        rom_memory[44660] = 3'b111;
        rom_memory[44661] = 3'b110;
        rom_memory[44662] = 3'b110;
        rom_memory[44663] = 3'b110;
        rom_memory[44664] = 3'b110;
        rom_memory[44665] = 3'b110;
        rom_memory[44666] = 3'b110;
        rom_memory[44667] = 3'b110;
        rom_memory[44668] = 3'b110;
        rom_memory[44669] = 3'b110;
        rom_memory[44670] = 3'b110;
        rom_memory[44671] = 3'b111;
        rom_memory[44672] = 3'b111;
        rom_memory[44673] = 3'b111;
        rom_memory[44674] = 3'b111;
        rom_memory[44675] = 3'b111;
        rom_memory[44676] = 3'b111;
        rom_memory[44677] = 3'b111;
        rom_memory[44678] = 3'b111;
        rom_memory[44679] = 3'b111;
        rom_memory[44680] = 3'b111;
        rom_memory[44681] = 3'b111;
        rom_memory[44682] = 3'b111;
        rom_memory[44683] = 3'b111;
        rom_memory[44684] = 3'b111;
        rom_memory[44685] = 3'b110;
        rom_memory[44686] = 3'b110;
        rom_memory[44687] = 3'b110;
        rom_memory[44688] = 3'b110;
        rom_memory[44689] = 3'b110;
        rom_memory[44690] = 3'b110;
        rom_memory[44691] = 3'b110;
        rom_memory[44692] = 3'b110;
        rom_memory[44693] = 3'b110;
        rom_memory[44694] = 3'b111;
        rom_memory[44695] = 3'b110;
        rom_memory[44696] = 3'b110;
        rom_memory[44697] = 3'b110;
        rom_memory[44698] = 3'b100;
        rom_memory[44699] = 3'b100;
        rom_memory[44700] = 3'b110;
        rom_memory[44701] = 3'b100;
        rom_memory[44702] = 3'b110;
        rom_memory[44703] = 3'b110;
        rom_memory[44704] = 3'b110;
        rom_memory[44705] = 3'b110;
        rom_memory[44706] = 3'b111;
        rom_memory[44707] = 3'b111;
        rom_memory[44708] = 3'b111;
        rom_memory[44709] = 3'b110;
        rom_memory[44710] = 3'b110;
        rom_memory[44711] = 3'b110;
        rom_memory[44712] = 3'b110;
        rom_memory[44713] = 3'b111;
        rom_memory[44714] = 3'b000;
        rom_memory[44715] = 3'b000;
        rom_memory[44716] = 3'b100;
        rom_memory[44717] = 3'b000;
        rom_memory[44718] = 3'b110;
        rom_memory[44719] = 3'b110;
        rom_memory[44720] = 3'b110;
        rom_memory[44721] = 3'b110;
        rom_memory[44722] = 3'b110;
        rom_memory[44723] = 3'b110;
        rom_memory[44724] = 3'b111;
        rom_memory[44725] = 3'b111;
        rom_memory[44726] = 3'b111;
        rom_memory[44727] = 3'b110;
        rom_memory[44728] = 3'b111;
        rom_memory[44729] = 3'b110;
        rom_memory[44730] = 3'b110;
        rom_memory[44731] = 3'b110;
        rom_memory[44732] = 3'b110;
        rom_memory[44733] = 3'b110;
        rom_memory[44734] = 3'b110;
        rom_memory[44735] = 3'b110;
        rom_memory[44736] = 3'b110;
        rom_memory[44737] = 3'b110;
        rom_memory[44738] = 3'b110;
        rom_memory[44739] = 3'b111;
        rom_memory[44740] = 3'b111;
        rom_memory[44741] = 3'b111;
        rom_memory[44742] = 3'b111;
        rom_memory[44743] = 3'b111;
        rom_memory[44744] = 3'b111;
        rom_memory[44745] = 3'b111;
        rom_memory[44746] = 3'b111;
        rom_memory[44747] = 3'b111;
        rom_memory[44748] = 3'b111;
        rom_memory[44749] = 3'b111;
        rom_memory[44750] = 3'b111;
        rom_memory[44751] = 3'b111;
        rom_memory[44752] = 3'b111;
        rom_memory[44753] = 3'b111;
        rom_memory[44754] = 3'b111;
        rom_memory[44755] = 3'b111;
        rom_memory[44756] = 3'b110;
        rom_memory[44757] = 3'b110;
        rom_memory[44758] = 3'b110;
        rom_memory[44759] = 3'b110;
        rom_memory[44760] = 3'b110;
        rom_memory[44761] = 3'b110;
        rom_memory[44762] = 3'b110;
        rom_memory[44763] = 3'b110;
        rom_memory[44764] = 3'b110;
        rom_memory[44765] = 3'b110;
        rom_memory[44766] = 3'b110;
        rom_memory[44767] = 3'b110;
        rom_memory[44768] = 3'b110;
        rom_memory[44769] = 3'b110;
        rom_memory[44770] = 3'b110;
        rom_memory[44771] = 3'b110;
        rom_memory[44772] = 3'b110;
        rom_memory[44773] = 3'b110;
        rom_memory[44774] = 3'b110;
        rom_memory[44775] = 3'b110;
        rom_memory[44776] = 3'b110;
        rom_memory[44777] = 3'b110;
        rom_memory[44778] = 3'b110;
        rom_memory[44779] = 3'b110;
        rom_memory[44780] = 3'b110;
        rom_memory[44781] = 3'b110;
        rom_memory[44782] = 3'b110;
        rom_memory[44783] = 3'b110;
        rom_memory[44784] = 3'b110;
        rom_memory[44785] = 3'b110;
        rom_memory[44786] = 3'b110;
        rom_memory[44787] = 3'b110;
        rom_memory[44788] = 3'b110;
        rom_memory[44789] = 3'b110;
        rom_memory[44790] = 3'b110;
        rom_memory[44791] = 3'b110;
        rom_memory[44792] = 3'b110;
        rom_memory[44793] = 3'b110;
        rom_memory[44794] = 3'b110;
        rom_memory[44795] = 3'b110;
        rom_memory[44796] = 3'b110;
        rom_memory[44797] = 3'b110;
        rom_memory[44798] = 3'b110;
        rom_memory[44799] = 3'b110;
        rom_memory[44800] = 3'b110;
        rom_memory[44801] = 3'b110;
        rom_memory[44802] = 3'b110;
        rom_memory[44803] = 3'b110;
        rom_memory[44804] = 3'b110;
        rom_memory[44805] = 3'b110;
        rom_memory[44806] = 3'b110;
        rom_memory[44807] = 3'b110;
        rom_memory[44808] = 3'b110;
        rom_memory[44809] = 3'b110;
        rom_memory[44810] = 3'b110;
        rom_memory[44811] = 3'b110;
        rom_memory[44812] = 3'b110;
        rom_memory[44813] = 3'b110;
        rom_memory[44814] = 3'b110;
        rom_memory[44815] = 3'b110;
        rom_memory[44816] = 3'b110;
        rom_memory[44817] = 3'b110;
        rom_memory[44818] = 3'b110;
        rom_memory[44819] = 3'b110;
        rom_memory[44820] = 3'b110;
        rom_memory[44821] = 3'b110;
        rom_memory[44822] = 3'b110;
        rom_memory[44823] = 3'b110;
        rom_memory[44824] = 3'b110;
        rom_memory[44825] = 3'b110;
        rom_memory[44826] = 3'b110;
        rom_memory[44827] = 3'b110;
        rom_memory[44828] = 3'b110;
        rom_memory[44829] = 3'b110;
        rom_memory[44830] = 3'b110;
        rom_memory[44831] = 3'b110;
        rom_memory[44832] = 3'b110;
        rom_memory[44833] = 3'b110;
        rom_memory[44834] = 3'b110;
        rom_memory[44835] = 3'b110;
        rom_memory[44836] = 3'b110;
        rom_memory[44837] = 3'b110;
        rom_memory[44838] = 3'b110;
        rom_memory[44839] = 3'b110;
        rom_memory[44840] = 3'b110;
        rom_memory[44841] = 3'b000;
        rom_memory[44842] = 3'b000;
        rom_memory[44843] = 3'b000;
        rom_memory[44844] = 3'b000;
        rom_memory[44845] = 3'b000;
        rom_memory[44846] = 3'b000;
        rom_memory[44847] = 3'b000;
        rom_memory[44848] = 3'b000;
        rom_memory[44849] = 3'b110;
        rom_memory[44850] = 3'b110;
        rom_memory[44851] = 3'b110;
        rom_memory[44852] = 3'b110;
        rom_memory[44853] = 3'b000;
        rom_memory[44854] = 3'b000;
        rom_memory[44855] = 3'b000;
        rom_memory[44856] = 3'b100;
        rom_memory[44857] = 3'b110;
        rom_memory[44858] = 3'b110;
        rom_memory[44859] = 3'b110;
        rom_memory[44860] = 3'b110;
        rom_memory[44861] = 3'b110;
        rom_memory[44862] = 3'b110;
        rom_memory[44863] = 3'b110;
        rom_memory[44864] = 3'b110;
        rom_memory[44865] = 3'b110;
        rom_memory[44866] = 3'b110;
        rom_memory[44867] = 3'b110;
        rom_memory[44868] = 3'b110;
        rom_memory[44869] = 3'b110;
        rom_memory[44870] = 3'b110;
        rom_memory[44871] = 3'b110;
        rom_memory[44872] = 3'b110;
        rom_memory[44873] = 3'b110;
        rom_memory[44874] = 3'b110;
        rom_memory[44875] = 3'b110;
        rom_memory[44876] = 3'b110;
        rom_memory[44877] = 3'b110;
        rom_memory[44878] = 3'b110;
        rom_memory[44879] = 3'b110;
        rom_memory[44880] = 3'b111;
        rom_memory[44881] = 3'b111;
        rom_memory[44882] = 3'b111;
        rom_memory[44883] = 3'b111;
        rom_memory[44884] = 3'b111;
        rom_memory[44885] = 3'b111;
        rom_memory[44886] = 3'b111;
        rom_memory[44887] = 3'b111;
        rom_memory[44888] = 3'b111;
        rom_memory[44889] = 3'b111;
        rom_memory[44890] = 3'b111;
        rom_memory[44891] = 3'b111;
        rom_memory[44892] = 3'b111;
        rom_memory[44893] = 3'b111;
        rom_memory[44894] = 3'b111;
        rom_memory[44895] = 3'b111;
        rom_memory[44896] = 3'b111;
        rom_memory[44897] = 3'b111;
        rom_memory[44898] = 3'b111;
        rom_memory[44899] = 3'b111;
        rom_memory[44900] = 3'b111;
        rom_memory[44901] = 3'b110;
        rom_memory[44902] = 3'b110;
        rom_memory[44903] = 3'b110;
        rom_memory[44904] = 3'b110;
        rom_memory[44905] = 3'b110;
        rom_memory[44906] = 3'b110;
        rom_memory[44907] = 3'b110;
        rom_memory[44908] = 3'b110;
        rom_memory[44909] = 3'b110;
        rom_memory[44910] = 3'b111;
        rom_memory[44911] = 3'b111;
        rom_memory[44912] = 3'b111;
        rom_memory[44913] = 3'b111;
        rom_memory[44914] = 3'b111;
        rom_memory[44915] = 3'b111;
        rom_memory[44916] = 3'b111;
        rom_memory[44917] = 3'b111;
        rom_memory[44918] = 3'b111;
        rom_memory[44919] = 3'b111;
        rom_memory[44920] = 3'b111;
        rom_memory[44921] = 3'b111;
        rom_memory[44922] = 3'b111;
        rom_memory[44923] = 3'b111;
        rom_memory[44924] = 3'b111;
        rom_memory[44925] = 3'b110;
        rom_memory[44926] = 3'b110;
        rom_memory[44927] = 3'b110;
        rom_memory[44928] = 3'b110;
        rom_memory[44929] = 3'b110;
        rom_memory[44930] = 3'b111;
        rom_memory[44931] = 3'b111;
        rom_memory[44932] = 3'b110;
        rom_memory[44933] = 3'b110;
        rom_memory[44934] = 3'b110;
        rom_memory[44935] = 3'b111;
        rom_memory[44936] = 3'b110;
        rom_memory[44937] = 3'b110;
        rom_memory[44938] = 3'b000;
        rom_memory[44939] = 3'b000;
        rom_memory[44940] = 3'b100;
        rom_memory[44941] = 3'b100;
        rom_memory[44942] = 3'b100;
        rom_memory[44943] = 3'b110;
        rom_memory[44944] = 3'b110;
        rom_memory[44945] = 3'b111;
        rom_memory[44946] = 3'b110;
        rom_memory[44947] = 3'b110;
        rom_memory[44948] = 3'b110;
        rom_memory[44949] = 3'b110;
        rom_memory[44950] = 3'b111;
        rom_memory[44951] = 3'b110;
        rom_memory[44952] = 3'b000;
        rom_memory[44953] = 3'b000;
        rom_memory[44954] = 3'b000;
        rom_memory[44955] = 3'b000;
        rom_memory[44956] = 3'b000;
        rom_memory[44957] = 3'b111;
        rom_memory[44958] = 3'b111;
        rom_memory[44959] = 3'b111;
        rom_memory[44960] = 3'b111;
        rom_memory[44961] = 3'b110;
        rom_memory[44962] = 3'b110;
        rom_memory[44963] = 3'b110;
        rom_memory[44964] = 3'b111;
        rom_memory[44965] = 3'b111;
        rom_memory[44966] = 3'b111;
        rom_memory[44967] = 3'b111;
        rom_memory[44968] = 3'b111;
        rom_memory[44969] = 3'b110;
        rom_memory[44970] = 3'b110;
        rom_memory[44971] = 3'b111;
        rom_memory[44972] = 3'b111;
        rom_memory[44973] = 3'b111;
        rom_memory[44974] = 3'b111;
        rom_memory[44975] = 3'b110;
        rom_memory[44976] = 3'b110;
        rom_memory[44977] = 3'b110;
        rom_memory[44978] = 3'b110;
        rom_memory[44979] = 3'b110;
        rom_memory[44980] = 3'b111;
        rom_memory[44981] = 3'b111;
        rom_memory[44982] = 3'b111;
        rom_memory[44983] = 3'b111;
        rom_memory[44984] = 3'b111;
        rom_memory[44985] = 3'b111;
        rom_memory[44986] = 3'b111;
        rom_memory[44987] = 3'b111;
        rom_memory[44988] = 3'b111;
        rom_memory[44989] = 3'b111;
        rom_memory[44990] = 3'b111;
        rom_memory[44991] = 3'b111;
        rom_memory[44992] = 3'b111;
        rom_memory[44993] = 3'b111;
        rom_memory[44994] = 3'b111;
        rom_memory[44995] = 3'b111;
        rom_memory[44996] = 3'b110;
        rom_memory[44997] = 3'b110;
        rom_memory[44998] = 3'b110;
        rom_memory[44999] = 3'b110;
        rom_memory[45000] = 3'b110;
        rom_memory[45001] = 3'b110;
        rom_memory[45002] = 3'b110;
        rom_memory[45003] = 3'b110;
        rom_memory[45004] = 3'b110;
        rom_memory[45005] = 3'b110;
        rom_memory[45006] = 3'b110;
        rom_memory[45007] = 3'b110;
        rom_memory[45008] = 3'b110;
        rom_memory[45009] = 3'b110;
        rom_memory[45010] = 3'b110;
        rom_memory[45011] = 3'b110;
        rom_memory[45012] = 3'b110;
        rom_memory[45013] = 3'b110;
        rom_memory[45014] = 3'b110;
        rom_memory[45015] = 3'b110;
        rom_memory[45016] = 3'b110;
        rom_memory[45017] = 3'b110;
        rom_memory[45018] = 3'b110;
        rom_memory[45019] = 3'b110;
        rom_memory[45020] = 3'b110;
        rom_memory[45021] = 3'b110;
        rom_memory[45022] = 3'b110;
        rom_memory[45023] = 3'b110;
        rom_memory[45024] = 3'b110;
        rom_memory[45025] = 3'b110;
        rom_memory[45026] = 3'b110;
        rom_memory[45027] = 3'b110;
        rom_memory[45028] = 3'b110;
        rom_memory[45029] = 3'b110;
        rom_memory[45030] = 3'b110;
        rom_memory[45031] = 3'b110;
        rom_memory[45032] = 3'b110;
        rom_memory[45033] = 3'b110;
        rom_memory[45034] = 3'b110;
        rom_memory[45035] = 3'b110;
        rom_memory[45036] = 3'b110;
        rom_memory[45037] = 3'b110;
        rom_memory[45038] = 3'b110;
        rom_memory[45039] = 3'b110;
        rom_memory[45040] = 3'b110;
        rom_memory[45041] = 3'b110;
        rom_memory[45042] = 3'b110;
        rom_memory[45043] = 3'b110;
        rom_memory[45044] = 3'b110;
        rom_memory[45045] = 3'b110;
        rom_memory[45046] = 3'b110;
        rom_memory[45047] = 3'b110;
        rom_memory[45048] = 3'b110;
        rom_memory[45049] = 3'b110;
        rom_memory[45050] = 3'b110;
        rom_memory[45051] = 3'b110;
        rom_memory[45052] = 3'b110;
        rom_memory[45053] = 3'b110;
        rom_memory[45054] = 3'b110;
        rom_memory[45055] = 3'b110;
        rom_memory[45056] = 3'b110;
        rom_memory[45057] = 3'b110;
        rom_memory[45058] = 3'b110;
        rom_memory[45059] = 3'b110;
        rom_memory[45060] = 3'b110;
        rom_memory[45061] = 3'b110;
        rom_memory[45062] = 3'b110;
        rom_memory[45063] = 3'b110;
        rom_memory[45064] = 3'b110;
        rom_memory[45065] = 3'b110;
        rom_memory[45066] = 3'b110;
        rom_memory[45067] = 3'b110;
        rom_memory[45068] = 3'b110;
        rom_memory[45069] = 3'b110;
        rom_memory[45070] = 3'b110;
        rom_memory[45071] = 3'b110;
        rom_memory[45072] = 3'b110;
        rom_memory[45073] = 3'b110;
        rom_memory[45074] = 3'b110;
        rom_memory[45075] = 3'b110;
        rom_memory[45076] = 3'b110;
        rom_memory[45077] = 3'b110;
        rom_memory[45078] = 3'b110;
        rom_memory[45079] = 3'b110;
        rom_memory[45080] = 3'b110;
        rom_memory[45081] = 3'b110;
        rom_memory[45082] = 3'b110;
        rom_memory[45083] = 3'b000;
        rom_memory[45084] = 3'b000;
        rom_memory[45085] = 3'b000;
        rom_memory[45086] = 3'b000;
        rom_memory[45087] = 3'b000;
        rom_memory[45088] = 3'b000;
        rom_memory[45089] = 3'b000;
        rom_memory[45090] = 3'b000;
        rom_memory[45091] = 3'b110;
        rom_memory[45092] = 3'b110;
        rom_memory[45093] = 3'b110;
        rom_memory[45094] = 3'b110;
        rom_memory[45095] = 3'b100;
        rom_memory[45096] = 3'b000;
        rom_memory[45097] = 3'b000;
        rom_memory[45098] = 3'b100;
        rom_memory[45099] = 3'b110;
        rom_memory[45100] = 3'b110;
        rom_memory[45101] = 3'b110;
        rom_memory[45102] = 3'b110;
        rom_memory[45103] = 3'b110;
        rom_memory[45104] = 3'b110;
        rom_memory[45105] = 3'b110;
        rom_memory[45106] = 3'b110;
        rom_memory[45107] = 3'b110;
        rom_memory[45108] = 3'b110;
        rom_memory[45109] = 3'b110;
        rom_memory[45110] = 3'b110;
        rom_memory[45111] = 3'b110;
        rom_memory[45112] = 3'b110;
        rom_memory[45113] = 3'b110;
        rom_memory[45114] = 3'b110;
        rom_memory[45115] = 3'b110;
        rom_memory[45116] = 3'b110;
        rom_memory[45117] = 3'b110;
        rom_memory[45118] = 3'b110;
        rom_memory[45119] = 3'b110;
        rom_memory[45120] = 3'b111;
        rom_memory[45121] = 3'b111;
        rom_memory[45122] = 3'b111;
        rom_memory[45123] = 3'b111;
        rom_memory[45124] = 3'b111;
        rom_memory[45125] = 3'b111;
        rom_memory[45126] = 3'b111;
        rom_memory[45127] = 3'b111;
        rom_memory[45128] = 3'b111;
        rom_memory[45129] = 3'b111;
        rom_memory[45130] = 3'b111;
        rom_memory[45131] = 3'b111;
        rom_memory[45132] = 3'b111;
        rom_memory[45133] = 3'b111;
        rom_memory[45134] = 3'b111;
        rom_memory[45135] = 3'b111;
        rom_memory[45136] = 3'b111;
        rom_memory[45137] = 3'b111;
        rom_memory[45138] = 3'b111;
        rom_memory[45139] = 3'b111;
        rom_memory[45140] = 3'b111;
        rom_memory[45141] = 3'b110;
        rom_memory[45142] = 3'b110;
        rom_memory[45143] = 3'b110;
        rom_memory[45144] = 3'b110;
        rom_memory[45145] = 3'b110;
        rom_memory[45146] = 3'b110;
        rom_memory[45147] = 3'b110;
        rom_memory[45148] = 3'b110;
        rom_memory[45149] = 3'b111;
        rom_memory[45150] = 3'b111;
        rom_memory[45151] = 3'b111;
        rom_memory[45152] = 3'b111;
        rom_memory[45153] = 3'b111;
        rom_memory[45154] = 3'b111;
        rom_memory[45155] = 3'b111;
        rom_memory[45156] = 3'b111;
        rom_memory[45157] = 3'b111;
        rom_memory[45158] = 3'b111;
        rom_memory[45159] = 3'b111;
        rom_memory[45160] = 3'b111;
        rom_memory[45161] = 3'b111;
        rom_memory[45162] = 3'b111;
        rom_memory[45163] = 3'b111;
        rom_memory[45164] = 3'b111;
        rom_memory[45165] = 3'b111;
        rom_memory[45166] = 3'b111;
        rom_memory[45167] = 3'b111;
        rom_memory[45168] = 3'b111;
        rom_memory[45169] = 3'b111;
        rom_memory[45170] = 3'b111;
        rom_memory[45171] = 3'b111;
        rom_memory[45172] = 3'b111;
        rom_memory[45173] = 3'b110;
        rom_memory[45174] = 3'b110;
        rom_memory[45175] = 3'b110;
        rom_memory[45176] = 3'b100;
        rom_memory[45177] = 3'b000;
        rom_memory[45178] = 3'b000;
        rom_memory[45179] = 3'b000;
        rom_memory[45180] = 3'b000;
        rom_memory[45181] = 3'b100;
        rom_memory[45182] = 3'b000;
        rom_memory[45183] = 3'b100;
        rom_memory[45184] = 3'b110;
        rom_memory[45185] = 3'b111;
        rom_memory[45186] = 3'b110;
        rom_memory[45187] = 3'b110;
        rom_memory[45188] = 3'b110;
        rom_memory[45189] = 3'b111;
        rom_memory[45190] = 3'b111;
        rom_memory[45191] = 3'b110;
        rom_memory[45192] = 3'b000;
        rom_memory[45193] = 3'b000;
        rom_memory[45194] = 3'b000;
        rom_memory[45195] = 3'b000;
        rom_memory[45196] = 3'b000;
        rom_memory[45197] = 3'b111;
        rom_memory[45198] = 3'b111;
        rom_memory[45199] = 3'b111;
        rom_memory[45200] = 3'b110;
        rom_memory[45201] = 3'b110;
        rom_memory[45202] = 3'b110;
        rom_memory[45203] = 3'b111;
        rom_memory[45204] = 3'b111;
        rom_memory[45205] = 3'b111;
        rom_memory[45206] = 3'b111;
        rom_memory[45207] = 3'b111;
        rom_memory[45208] = 3'b111;
        rom_memory[45209] = 3'b111;
        rom_memory[45210] = 3'b111;
        rom_memory[45211] = 3'b111;
        rom_memory[45212] = 3'b111;
        rom_memory[45213] = 3'b111;
        rom_memory[45214] = 3'b111;
        rom_memory[45215] = 3'b111;
        rom_memory[45216] = 3'b111;
        rom_memory[45217] = 3'b110;
        rom_memory[45218] = 3'b110;
        rom_memory[45219] = 3'b110;
        rom_memory[45220] = 3'b110;
        rom_memory[45221] = 3'b110;
        rom_memory[45222] = 3'b111;
        rom_memory[45223] = 3'b111;
        rom_memory[45224] = 3'b111;
        rom_memory[45225] = 3'b111;
        rom_memory[45226] = 3'b111;
        rom_memory[45227] = 3'b111;
        rom_memory[45228] = 3'b111;
        rom_memory[45229] = 3'b111;
        rom_memory[45230] = 3'b111;
        rom_memory[45231] = 3'b111;
        rom_memory[45232] = 3'b111;
        rom_memory[45233] = 3'b111;
        rom_memory[45234] = 3'b111;
        rom_memory[45235] = 3'b111;
        rom_memory[45236] = 3'b110;
        rom_memory[45237] = 3'b110;
        rom_memory[45238] = 3'b110;
        rom_memory[45239] = 3'b110;
        rom_memory[45240] = 3'b110;
        rom_memory[45241] = 3'b110;
        rom_memory[45242] = 3'b110;
        rom_memory[45243] = 3'b110;
        rom_memory[45244] = 3'b110;
        rom_memory[45245] = 3'b110;
        rom_memory[45246] = 3'b110;
        rom_memory[45247] = 3'b110;
        rom_memory[45248] = 3'b110;
        rom_memory[45249] = 3'b110;
        rom_memory[45250] = 3'b110;
        rom_memory[45251] = 3'b110;
        rom_memory[45252] = 3'b110;
        rom_memory[45253] = 3'b110;
        rom_memory[45254] = 3'b110;
        rom_memory[45255] = 3'b110;
        rom_memory[45256] = 3'b110;
        rom_memory[45257] = 3'b110;
        rom_memory[45258] = 3'b110;
        rom_memory[45259] = 3'b110;
        rom_memory[45260] = 3'b110;
        rom_memory[45261] = 3'b110;
        rom_memory[45262] = 3'b110;
        rom_memory[45263] = 3'b110;
        rom_memory[45264] = 3'b110;
        rom_memory[45265] = 3'b110;
        rom_memory[45266] = 3'b110;
        rom_memory[45267] = 3'b110;
        rom_memory[45268] = 3'b110;
        rom_memory[45269] = 3'b110;
        rom_memory[45270] = 3'b110;
        rom_memory[45271] = 3'b110;
        rom_memory[45272] = 3'b110;
        rom_memory[45273] = 3'b110;
        rom_memory[45274] = 3'b110;
        rom_memory[45275] = 3'b110;
        rom_memory[45276] = 3'b110;
        rom_memory[45277] = 3'b110;
        rom_memory[45278] = 3'b110;
        rom_memory[45279] = 3'b110;
        rom_memory[45280] = 3'b110;
        rom_memory[45281] = 3'b110;
        rom_memory[45282] = 3'b110;
        rom_memory[45283] = 3'b110;
        rom_memory[45284] = 3'b110;
        rom_memory[45285] = 3'b110;
        rom_memory[45286] = 3'b110;
        rom_memory[45287] = 3'b110;
        rom_memory[45288] = 3'b110;
        rom_memory[45289] = 3'b110;
        rom_memory[45290] = 3'b110;
        rom_memory[45291] = 3'b110;
        rom_memory[45292] = 3'b110;
        rom_memory[45293] = 3'b110;
        rom_memory[45294] = 3'b110;
        rom_memory[45295] = 3'b110;
        rom_memory[45296] = 3'b110;
        rom_memory[45297] = 3'b110;
        rom_memory[45298] = 3'b110;
        rom_memory[45299] = 3'b110;
        rom_memory[45300] = 3'b110;
        rom_memory[45301] = 3'b110;
        rom_memory[45302] = 3'b110;
        rom_memory[45303] = 3'b110;
        rom_memory[45304] = 3'b110;
        rom_memory[45305] = 3'b110;
        rom_memory[45306] = 3'b110;
        rom_memory[45307] = 3'b110;
        rom_memory[45308] = 3'b110;
        rom_memory[45309] = 3'b110;
        rom_memory[45310] = 3'b110;
        rom_memory[45311] = 3'b110;
        rom_memory[45312] = 3'b110;
        rom_memory[45313] = 3'b110;
        rom_memory[45314] = 3'b110;
        rom_memory[45315] = 3'b110;
        rom_memory[45316] = 3'b110;
        rom_memory[45317] = 3'b110;
        rom_memory[45318] = 3'b110;
        rom_memory[45319] = 3'b110;
        rom_memory[45320] = 3'b110;
        rom_memory[45321] = 3'b110;
        rom_memory[45322] = 3'b110;
        rom_memory[45323] = 3'b110;
        rom_memory[45324] = 3'b100;
        rom_memory[45325] = 3'b000;
        rom_memory[45326] = 3'b000;
        rom_memory[45327] = 3'b000;
        rom_memory[45328] = 3'b000;
        rom_memory[45329] = 3'b000;
        rom_memory[45330] = 3'b000;
        rom_memory[45331] = 3'b000;
        rom_memory[45332] = 3'b100;
        rom_memory[45333] = 3'b110;
        rom_memory[45334] = 3'b110;
        rom_memory[45335] = 3'b110;
        rom_memory[45336] = 3'b110;
        rom_memory[45337] = 3'b110;
        rom_memory[45338] = 3'b100;
        rom_memory[45339] = 3'b000;
        rom_memory[45340] = 3'b100;
        rom_memory[45341] = 3'b110;
        rom_memory[45342] = 3'b110;
        rom_memory[45343] = 3'b110;
        rom_memory[45344] = 3'b110;
        rom_memory[45345] = 3'b110;
        rom_memory[45346] = 3'b110;
        rom_memory[45347] = 3'b110;
        rom_memory[45348] = 3'b110;
        rom_memory[45349] = 3'b110;
        rom_memory[45350] = 3'b110;
        rom_memory[45351] = 3'b110;
        rom_memory[45352] = 3'b110;
        rom_memory[45353] = 3'b110;
        rom_memory[45354] = 3'b110;
        rom_memory[45355] = 3'b110;
        rom_memory[45356] = 3'b110;
        rom_memory[45357] = 3'b110;
        rom_memory[45358] = 3'b110;
        rom_memory[45359] = 3'b110;
        rom_memory[45360] = 3'b111;
        rom_memory[45361] = 3'b111;
        rom_memory[45362] = 3'b111;
        rom_memory[45363] = 3'b111;
        rom_memory[45364] = 3'b111;
        rom_memory[45365] = 3'b111;
        rom_memory[45366] = 3'b111;
        rom_memory[45367] = 3'b111;
        rom_memory[45368] = 3'b111;
        rom_memory[45369] = 3'b111;
        rom_memory[45370] = 3'b111;
        rom_memory[45371] = 3'b111;
        rom_memory[45372] = 3'b111;
        rom_memory[45373] = 3'b111;
        rom_memory[45374] = 3'b111;
        rom_memory[45375] = 3'b111;
        rom_memory[45376] = 3'b111;
        rom_memory[45377] = 3'b111;
        rom_memory[45378] = 3'b111;
        rom_memory[45379] = 3'b111;
        rom_memory[45380] = 3'b110;
        rom_memory[45381] = 3'b110;
        rom_memory[45382] = 3'b110;
        rom_memory[45383] = 3'b110;
        rom_memory[45384] = 3'b110;
        rom_memory[45385] = 3'b110;
        rom_memory[45386] = 3'b110;
        rom_memory[45387] = 3'b110;
        rom_memory[45388] = 3'b110;
        rom_memory[45389] = 3'b110;
        rom_memory[45390] = 3'b111;
        rom_memory[45391] = 3'b111;
        rom_memory[45392] = 3'b111;
        rom_memory[45393] = 3'b111;
        rom_memory[45394] = 3'b111;
        rom_memory[45395] = 3'b111;
        rom_memory[45396] = 3'b111;
        rom_memory[45397] = 3'b111;
        rom_memory[45398] = 3'b111;
        rom_memory[45399] = 3'b111;
        rom_memory[45400] = 3'b111;
        rom_memory[45401] = 3'b111;
        rom_memory[45402] = 3'b111;
        rom_memory[45403] = 3'b111;
        rom_memory[45404] = 3'b111;
        rom_memory[45405] = 3'b111;
        rom_memory[45406] = 3'b111;
        rom_memory[45407] = 3'b111;
        rom_memory[45408] = 3'b111;
        rom_memory[45409] = 3'b111;
        rom_memory[45410] = 3'b111;
        rom_memory[45411] = 3'b111;
        rom_memory[45412] = 3'b110;
        rom_memory[45413] = 3'b110;
        rom_memory[45414] = 3'b110;
        rom_memory[45415] = 3'b110;
        rom_memory[45416] = 3'b110;
        rom_memory[45417] = 3'b100;
        rom_memory[45418] = 3'b100;
        rom_memory[45419] = 3'b000;
        rom_memory[45420] = 3'b000;
        rom_memory[45421] = 3'b000;
        rom_memory[45422] = 3'b100;
        rom_memory[45423] = 3'b100;
        rom_memory[45424] = 3'b111;
        rom_memory[45425] = 3'b111;
        rom_memory[45426] = 3'b111;
        rom_memory[45427] = 3'b110;
        rom_memory[45428] = 3'b110;
        rom_memory[45429] = 3'b111;
        rom_memory[45430] = 3'b110;
        rom_memory[45431] = 3'b000;
        rom_memory[45432] = 3'b000;
        rom_memory[45433] = 3'b000;
        rom_memory[45434] = 3'b000;
        rom_memory[45435] = 3'b000;
        rom_memory[45436] = 3'b111;
        rom_memory[45437] = 3'b111;
        rom_memory[45438] = 3'b111;
        rom_memory[45439] = 3'b110;
        rom_memory[45440] = 3'b110;
        rom_memory[45441] = 3'b110;
        rom_memory[45442] = 3'b110;
        rom_memory[45443] = 3'b111;
        rom_memory[45444] = 3'b111;
        rom_memory[45445] = 3'b111;
        rom_memory[45446] = 3'b111;
        rom_memory[45447] = 3'b111;
        rom_memory[45448] = 3'b111;
        rom_memory[45449] = 3'b111;
        rom_memory[45450] = 3'b111;
        rom_memory[45451] = 3'b111;
        rom_memory[45452] = 3'b111;
        rom_memory[45453] = 3'b111;
        rom_memory[45454] = 3'b111;
        rom_memory[45455] = 3'b111;
        rom_memory[45456] = 3'b110;
        rom_memory[45457] = 3'b110;
        rom_memory[45458] = 3'b110;
        rom_memory[45459] = 3'b110;
        rom_memory[45460] = 3'b110;
        rom_memory[45461] = 3'b110;
        rom_memory[45462] = 3'b110;
        rom_memory[45463] = 3'b111;
        rom_memory[45464] = 3'b111;
        rom_memory[45465] = 3'b111;
        rom_memory[45466] = 3'b111;
        rom_memory[45467] = 3'b111;
        rom_memory[45468] = 3'b111;
        rom_memory[45469] = 3'b111;
        rom_memory[45470] = 3'b111;
        rom_memory[45471] = 3'b111;
        rom_memory[45472] = 3'b111;
        rom_memory[45473] = 3'b111;
        rom_memory[45474] = 3'b111;
        rom_memory[45475] = 3'b111;
        rom_memory[45476] = 3'b110;
        rom_memory[45477] = 3'b110;
        rom_memory[45478] = 3'b110;
        rom_memory[45479] = 3'b110;
        rom_memory[45480] = 3'b110;
        rom_memory[45481] = 3'b110;
        rom_memory[45482] = 3'b110;
        rom_memory[45483] = 3'b110;
        rom_memory[45484] = 3'b110;
        rom_memory[45485] = 3'b110;
        rom_memory[45486] = 3'b110;
        rom_memory[45487] = 3'b110;
        rom_memory[45488] = 3'b110;
        rom_memory[45489] = 3'b110;
        rom_memory[45490] = 3'b110;
        rom_memory[45491] = 3'b110;
        rom_memory[45492] = 3'b110;
        rom_memory[45493] = 3'b110;
        rom_memory[45494] = 3'b110;
        rom_memory[45495] = 3'b110;
        rom_memory[45496] = 3'b110;
        rom_memory[45497] = 3'b110;
        rom_memory[45498] = 3'b110;
        rom_memory[45499] = 3'b110;
        rom_memory[45500] = 3'b110;
        rom_memory[45501] = 3'b110;
        rom_memory[45502] = 3'b110;
        rom_memory[45503] = 3'b110;
        rom_memory[45504] = 3'b110;
        rom_memory[45505] = 3'b110;
        rom_memory[45506] = 3'b110;
        rom_memory[45507] = 3'b110;
        rom_memory[45508] = 3'b110;
        rom_memory[45509] = 3'b110;
        rom_memory[45510] = 3'b110;
        rom_memory[45511] = 3'b110;
        rom_memory[45512] = 3'b110;
        rom_memory[45513] = 3'b110;
        rom_memory[45514] = 3'b110;
        rom_memory[45515] = 3'b110;
        rom_memory[45516] = 3'b110;
        rom_memory[45517] = 3'b110;
        rom_memory[45518] = 3'b110;
        rom_memory[45519] = 3'b110;
        rom_memory[45520] = 3'b110;
        rom_memory[45521] = 3'b110;
        rom_memory[45522] = 3'b110;
        rom_memory[45523] = 3'b110;
        rom_memory[45524] = 3'b110;
        rom_memory[45525] = 3'b110;
        rom_memory[45526] = 3'b110;
        rom_memory[45527] = 3'b110;
        rom_memory[45528] = 3'b110;
        rom_memory[45529] = 3'b110;
        rom_memory[45530] = 3'b110;
        rom_memory[45531] = 3'b110;
        rom_memory[45532] = 3'b110;
        rom_memory[45533] = 3'b110;
        rom_memory[45534] = 3'b110;
        rom_memory[45535] = 3'b110;
        rom_memory[45536] = 3'b110;
        rom_memory[45537] = 3'b110;
        rom_memory[45538] = 3'b110;
        rom_memory[45539] = 3'b110;
        rom_memory[45540] = 3'b110;
        rom_memory[45541] = 3'b110;
        rom_memory[45542] = 3'b110;
        rom_memory[45543] = 3'b110;
        rom_memory[45544] = 3'b110;
        rom_memory[45545] = 3'b110;
        rom_memory[45546] = 3'b110;
        rom_memory[45547] = 3'b110;
        rom_memory[45548] = 3'b110;
        rom_memory[45549] = 3'b110;
        rom_memory[45550] = 3'b110;
        rom_memory[45551] = 3'b110;
        rom_memory[45552] = 3'b110;
        rom_memory[45553] = 3'b110;
        rom_memory[45554] = 3'b110;
        rom_memory[45555] = 3'b110;
        rom_memory[45556] = 3'b110;
        rom_memory[45557] = 3'b110;
        rom_memory[45558] = 3'b110;
        rom_memory[45559] = 3'b110;
        rom_memory[45560] = 3'b110;
        rom_memory[45561] = 3'b110;
        rom_memory[45562] = 3'b110;
        rom_memory[45563] = 3'b110;
        rom_memory[45564] = 3'b110;
        rom_memory[45565] = 3'b110;
        rom_memory[45566] = 3'b100;
        rom_memory[45567] = 3'b000;
        rom_memory[45568] = 3'b000;
        rom_memory[45569] = 3'b000;
        rom_memory[45570] = 3'b000;
        rom_memory[45571] = 3'b000;
        rom_memory[45572] = 3'b000;
        rom_memory[45573] = 3'b000;
        rom_memory[45574] = 3'b110;
        rom_memory[45575] = 3'b110;
        rom_memory[45576] = 3'b110;
        rom_memory[45577] = 3'b110;
        rom_memory[45578] = 3'b110;
        rom_memory[45579] = 3'b110;
        rom_memory[45580] = 3'b100;
        rom_memory[45581] = 3'b000;
        rom_memory[45582] = 3'b100;
        rom_memory[45583] = 3'b110;
        rom_memory[45584] = 3'b110;
        rom_memory[45585] = 3'b110;
        rom_memory[45586] = 3'b110;
        rom_memory[45587] = 3'b110;
        rom_memory[45588] = 3'b110;
        rom_memory[45589] = 3'b110;
        rom_memory[45590] = 3'b110;
        rom_memory[45591] = 3'b110;
        rom_memory[45592] = 3'b110;
        rom_memory[45593] = 3'b110;
        rom_memory[45594] = 3'b110;
        rom_memory[45595] = 3'b110;
        rom_memory[45596] = 3'b110;
        rom_memory[45597] = 3'b110;
        rom_memory[45598] = 3'b110;
        rom_memory[45599] = 3'b110;
        rom_memory[45600] = 3'b111;
        rom_memory[45601] = 3'b111;
        rom_memory[45602] = 3'b111;
        rom_memory[45603] = 3'b111;
        rom_memory[45604] = 3'b111;
        rom_memory[45605] = 3'b111;
        rom_memory[45606] = 3'b111;
        rom_memory[45607] = 3'b111;
        rom_memory[45608] = 3'b111;
        rom_memory[45609] = 3'b111;
        rom_memory[45610] = 3'b111;
        rom_memory[45611] = 3'b111;
        rom_memory[45612] = 3'b111;
        rom_memory[45613] = 3'b111;
        rom_memory[45614] = 3'b111;
        rom_memory[45615] = 3'b111;
        rom_memory[45616] = 3'b111;
        rom_memory[45617] = 3'b111;
        rom_memory[45618] = 3'b111;
        rom_memory[45619] = 3'b111;
        rom_memory[45620] = 3'b110;
        rom_memory[45621] = 3'b110;
        rom_memory[45622] = 3'b110;
        rom_memory[45623] = 3'b110;
        rom_memory[45624] = 3'b110;
        rom_memory[45625] = 3'b110;
        rom_memory[45626] = 3'b110;
        rom_memory[45627] = 3'b110;
        rom_memory[45628] = 3'b110;
        rom_memory[45629] = 3'b110;
        rom_memory[45630] = 3'b111;
        rom_memory[45631] = 3'b111;
        rom_memory[45632] = 3'b111;
        rom_memory[45633] = 3'b111;
        rom_memory[45634] = 3'b111;
        rom_memory[45635] = 3'b111;
        rom_memory[45636] = 3'b111;
        rom_memory[45637] = 3'b111;
        rom_memory[45638] = 3'b111;
        rom_memory[45639] = 3'b111;
        rom_memory[45640] = 3'b111;
        rom_memory[45641] = 3'b111;
        rom_memory[45642] = 3'b111;
        rom_memory[45643] = 3'b111;
        rom_memory[45644] = 3'b111;
        rom_memory[45645] = 3'b111;
        rom_memory[45646] = 3'b111;
        rom_memory[45647] = 3'b111;
        rom_memory[45648] = 3'b111;
        rom_memory[45649] = 3'b111;
        rom_memory[45650] = 3'b111;
        rom_memory[45651] = 3'b111;
        rom_memory[45652] = 3'b110;
        rom_memory[45653] = 3'b110;
        rom_memory[45654] = 3'b110;
        rom_memory[45655] = 3'b110;
        rom_memory[45656] = 3'b110;
        rom_memory[45657] = 3'b100;
        rom_memory[45658] = 3'b100;
        rom_memory[45659] = 3'b100;
        rom_memory[45660] = 3'b000;
        rom_memory[45661] = 3'b000;
        rom_memory[45662] = 3'b000;
        rom_memory[45663] = 3'b100;
        rom_memory[45664] = 3'b111;
        rom_memory[45665] = 3'b111;
        rom_memory[45666] = 3'b111;
        rom_memory[45667] = 3'b110;
        rom_memory[45668] = 3'b110;
        rom_memory[45669] = 3'b111;
        rom_memory[45670] = 3'b110;
        rom_memory[45671] = 3'b000;
        rom_memory[45672] = 3'b110;
        rom_memory[45673] = 3'b000;
        rom_memory[45674] = 3'b000;
        rom_memory[45675] = 3'b000;
        rom_memory[45676] = 3'b111;
        rom_memory[45677] = 3'b111;
        rom_memory[45678] = 3'b111;
        rom_memory[45679] = 3'b110;
        rom_memory[45680] = 3'b110;
        rom_memory[45681] = 3'b111;
        rom_memory[45682] = 3'b111;
        rom_memory[45683] = 3'b111;
        rom_memory[45684] = 3'b111;
        rom_memory[45685] = 3'b111;
        rom_memory[45686] = 3'b111;
        rom_memory[45687] = 3'b111;
        rom_memory[45688] = 3'b111;
        rom_memory[45689] = 3'b111;
        rom_memory[45690] = 3'b111;
        rom_memory[45691] = 3'b111;
        rom_memory[45692] = 3'b111;
        rom_memory[45693] = 3'b111;
        rom_memory[45694] = 3'b111;
        rom_memory[45695] = 3'b110;
        rom_memory[45696] = 3'b110;
        rom_memory[45697] = 3'b110;
        rom_memory[45698] = 3'b110;
        rom_memory[45699] = 3'b110;
        rom_memory[45700] = 3'b110;
        rom_memory[45701] = 3'b100;
        rom_memory[45702] = 3'b100;
        rom_memory[45703] = 3'b110;
        rom_memory[45704] = 3'b111;
        rom_memory[45705] = 3'b111;
        rom_memory[45706] = 3'b111;
        rom_memory[45707] = 3'b111;
        rom_memory[45708] = 3'b111;
        rom_memory[45709] = 3'b111;
        rom_memory[45710] = 3'b111;
        rom_memory[45711] = 3'b111;
        rom_memory[45712] = 3'b111;
        rom_memory[45713] = 3'b111;
        rom_memory[45714] = 3'b111;
        rom_memory[45715] = 3'b111;
        rom_memory[45716] = 3'b110;
        rom_memory[45717] = 3'b110;
        rom_memory[45718] = 3'b110;
        rom_memory[45719] = 3'b110;
        rom_memory[45720] = 3'b110;
        rom_memory[45721] = 3'b110;
        rom_memory[45722] = 3'b110;
        rom_memory[45723] = 3'b110;
        rom_memory[45724] = 3'b110;
        rom_memory[45725] = 3'b110;
        rom_memory[45726] = 3'b110;
        rom_memory[45727] = 3'b110;
        rom_memory[45728] = 3'b110;
        rom_memory[45729] = 3'b110;
        rom_memory[45730] = 3'b110;
        rom_memory[45731] = 3'b110;
        rom_memory[45732] = 3'b110;
        rom_memory[45733] = 3'b110;
        rom_memory[45734] = 3'b110;
        rom_memory[45735] = 3'b110;
        rom_memory[45736] = 3'b110;
        rom_memory[45737] = 3'b110;
        rom_memory[45738] = 3'b110;
        rom_memory[45739] = 3'b110;
        rom_memory[45740] = 3'b110;
        rom_memory[45741] = 3'b110;
        rom_memory[45742] = 3'b110;
        rom_memory[45743] = 3'b110;
        rom_memory[45744] = 3'b110;
        rom_memory[45745] = 3'b110;
        rom_memory[45746] = 3'b110;
        rom_memory[45747] = 3'b110;
        rom_memory[45748] = 3'b110;
        rom_memory[45749] = 3'b110;
        rom_memory[45750] = 3'b110;
        rom_memory[45751] = 3'b110;
        rom_memory[45752] = 3'b110;
        rom_memory[45753] = 3'b110;
        rom_memory[45754] = 3'b110;
        rom_memory[45755] = 3'b110;
        rom_memory[45756] = 3'b110;
        rom_memory[45757] = 3'b110;
        rom_memory[45758] = 3'b110;
        rom_memory[45759] = 3'b110;
        rom_memory[45760] = 3'b110;
        rom_memory[45761] = 3'b110;
        rom_memory[45762] = 3'b110;
        rom_memory[45763] = 3'b110;
        rom_memory[45764] = 3'b110;
        rom_memory[45765] = 3'b110;
        rom_memory[45766] = 3'b110;
        rom_memory[45767] = 3'b110;
        rom_memory[45768] = 3'b110;
        rom_memory[45769] = 3'b110;
        rom_memory[45770] = 3'b110;
        rom_memory[45771] = 3'b110;
        rom_memory[45772] = 3'b110;
        rom_memory[45773] = 3'b110;
        rom_memory[45774] = 3'b110;
        rom_memory[45775] = 3'b110;
        rom_memory[45776] = 3'b110;
        rom_memory[45777] = 3'b110;
        rom_memory[45778] = 3'b110;
        rom_memory[45779] = 3'b110;
        rom_memory[45780] = 3'b110;
        rom_memory[45781] = 3'b110;
        rom_memory[45782] = 3'b110;
        rom_memory[45783] = 3'b110;
        rom_memory[45784] = 3'b110;
        rom_memory[45785] = 3'b110;
        rom_memory[45786] = 3'b110;
        rom_memory[45787] = 3'b110;
        rom_memory[45788] = 3'b110;
        rom_memory[45789] = 3'b110;
        rom_memory[45790] = 3'b110;
        rom_memory[45791] = 3'b110;
        rom_memory[45792] = 3'b110;
        rom_memory[45793] = 3'b110;
        rom_memory[45794] = 3'b110;
        rom_memory[45795] = 3'b110;
        rom_memory[45796] = 3'b110;
        rom_memory[45797] = 3'b110;
        rom_memory[45798] = 3'b110;
        rom_memory[45799] = 3'b110;
        rom_memory[45800] = 3'b110;
        rom_memory[45801] = 3'b110;
        rom_memory[45802] = 3'b110;
        rom_memory[45803] = 3'b110;
        rom_memory[45804] = 3'b110;
        rom_memory[45805] = 3'b110;
        rom_memory[45806] = 3'b110;
        rom_memory[45807] = 3'b110;
        rom_memory[45808] = 3'b100;
        rom_memory[45809] = 3'b000;
        rom_memory[45810] = 3'b000;
        rom_memory[45811] = 3'b000;
        rom_memory[45812] = 3'b000;
        rom_memory[45813] = 3'b000;
        rom_memory[45814] = 3'b000;
        rom_memory[45815] = 3'b000;
        rom_memory[45816] = 3'b110;
        rom_memory[45817] = 3'b110;
        rom_memory[45818] = 3'b110;
        rom_memory[45819] = 3'b110;
        rom_memory[45820] = 3'b110;
        rom_memory[45821] = 3'b110;
        rom_memory[45822] = 3'b110;
        rom_memory[45823] = 3'b100;
        rom_memory[45824] = 3'b100;
        rom_memory[45825] = 3'b110;
        rom_memory[45826] = 3'b110;
        rom_memory[45827] = 3'b110;
        rom_memory[45828] = 3'b110;
        rom_memory[45829] = 3'b110;
        rom_memory[45830] = 3'b110;
        rom_memory[45831] = 3'b110;
        rom_memory[45832] = 3'b110;
        rom_memory[45833] = 3'b110;
        rom_memory[45834] = 3'b110;
        rom_memory[45835] = 3'b110;
        rom_memory[45836] = 3'b110;
        rom_memory[45837] = 3'b110;
        rom_memory[45838] = 3'b110;
        rom_memory[45839] = 3'b110;
        rom_memory[45840] = 3'b110;
        rom_memory[45841] = 3'b111;
        rom_memory[45842] = 3'b111;
        rom_memory[45843] = 3'b111;
        rom_memory[45844] = 3'b111;
        rom_memory[45845] = 3'b111;
        rom_memory[45846] = 3'b111;
        rom_memory[45847] = 3'b111;
        rom_memory[45848] = 3'b111;
        rom_memory[45849] = 3'b111;
        rom_memory[45850] = 3'b111;
        rom_memory[45851] = 3'b111;
        rom_memory[45852] = 3'b111;
        rom_memory[45853] = 3'b111;
        rom_memory[45854] = 3'b111;
        rom_memory[45855] = 3'b111;
        rom_memory[45856] = 3'b111;
        rom_memory[45857] = 3'b111;
        rom_memory[45858] = 3'b111;
        rom_memory[45859] = 3'b111;
        rom_memory[45860] = 3'b111;
        rom_memory[45861] = 3'b110;
        rom_memory[45862] = 3'b110;
        rom_memory[45863] = 3'b110;
        rom_memory[45864] = 3'b110;
        rom_memory[45865] = 3'b110;
        rom_memory[45866] = 3'b110;
        rom_memory[45867] = 3'b110;
        rom_memory[45868] = 3'b110;
        rom_memory[45869] = 3'b110;
        rom_memory[45870] = 3'b111;
        rom_memory[45871] = 3'b111;
        rom_memory[45872] = 3'b111;
        rom_memory[45873] = 3'b111;
        rom_memory[45874] = 3'b111;
        rom_memory[45875] = 3'b111;
        rom_memory[45876] = 3'b111;
        rom_memory[45877] = 3'b111;
        rom_memory[45878] = 3'b111;
        rom_memory[45879] = 3'b111;
        rom_memory[45880] = 3'b111;
        rom_memory[45881] = 3'b111;
        rom_memory[45882] = 3'b111;
        rom_memory[45883] = 3'b111;
        rom_memory[45884] = 3'b111;
        rom_memory[45885] = 3'b111;
        rom_memory[45886] = 3'b111;
        rom_memory[45887] = 3'b111;
        rom_memory[45888] = 3'b111;
        rom_memory[45889] = 3'b111;
        rom_memory[45890] = 3'b111;
        rom_memory[45891] = 3'b110;
        rom_memory[45892] = 3'b110;
        rom_memory[45893] = 3'b110;
        rom_memory[45894] = 3'b110;
        rom_memory[45895] = 3'b111;
        rom_memory[45896] = 3'b110;
        rom_memory[45897] = 3'b100;
        rom_memory[45898] = 3'b100;
        rom_memory[45899] = 3'b100;
        rom_memory[45900] = 3'b100;
        rom_memory[45901] = 3'b000;
        rom_memory[45902] = 3'b000;
        rom_memory[45903] = 3'b100;
        rom_memory[45904] = 3'b100;
        rom_memory[45905] = 3'b111;
        rom_memory[45906] = 3'b111;
        rom_memory[45907] = 3'b111;
        rom_memory[45908] = 3'b111;
        rom_memory[45909] = 3'b111;
        rom_memory[45910] = 3'b110;
        rom_memory[45911] = 3'b100;
        rom_memory[45912] = 3'b100;
        rom_memory[45913] = 3'b100;
        rom_memory[45914] = 3'b000;
        rom_memory[45915] = 3'b110;
        rom_memory[45916] = 3'b111;
        rom_memory[45917] = 3'b111;
        rom_memory[45918] = 3'b111;
        rom_memory[45919] = 3'b111;
        rom_memory[45920] = 3'b111;
        rom_memory[45921] = 3'b111;
        rom_memory[45922] = 3'b111;
        rom_memory[45923] = 3'b111;
        rom_memory[45924] = 3'b111;
        rom_memory[45925] = 3'b111;
        rom_memory[45926] = 3'b111;
        rom_memory[45927] = 3'b111;
        rom_memory[45928] = 3'b111;
        rom_memory[45929] = 3'b111;
        rom_memory[45930] = 3'b111;
        rom_memory[45931] = 3'b111;
        rom_memory[45932] = 3'b111;
        rom_memory[45933] = 3'b111;
        rom_memory[45934] = 3'b110;
        rom_memory[45935] = 3'b110;
        rom_memory[45936] = 3'b110;
        rom_memory[45937] = 3'b110;
        rom_memory[45938] = 3'b110;
        rom_memory[45939] = 3'b110;
        rom_memory[45940] = 3'b110;
        rom_memory[45941] = 3'b110;
        rom_memory[45942] = 3'b110;
        rom_memory[45943] = 3'b110;
        rom_memory[45944] = 3'b111;
        rom_memory[45945] = 3'b111;
        rom_memory[45946] = 3'b111;
        rom_memory[45947] = 3'b111;
        rom_memory[45948] = 3'b111;
        rom_memory[45949] = 3'b111;
        rom_memory[45950] = 3'b111;
        rom_memory[45951] = 3'b111;
        rom_memory[45952] = 3'b111;
        rom_memory[45953] = 3'b111;
        rom_memory[45954] = 3'b111;
        rom_memory[45955] = 3'b111;
        rom_memory[45956] = 3'b110;
        rom_memory[45957] = 3'b110;
        rom_memory[45958] = 3'b110;
        rom_memory[45959] = 3'b110;
        rom_memory[45960] = 3'b110;
        rom_memory[45961] = 3'b110;
        rom_memory[45962] = 3'b110;
        rom_memory[45963] = 3'b110;
        rom_memory[45964] = 3'b110;
        rom_memory[45965] = 3'b110;
        rom_memory[45966] = 3'b110;
        rom_memory[45967] = 3'b110;
        rom_memory[45968] = 3'b110;
        rom_memory[45969] = 3'b110;
        rom_memory[45970] = 3'b110;
        rom_memory[45971] = 3'b110;
        rom_memory[45972] = 3'b110;
        rom_memory[45973] = 3'b110;
        rom_memory[45974] = 3'b110;
        rom_memory[45975] = 3'b110;
        rom_memory[45976] = 3'b110;
        rom_memory[45977] = 3'b110;
        rom_memory[45978] = 3'b110;
        rom_memory[45979] = 3'b110;
        rom_memory[45980] = 3'b110;
        rom_memory[45981] = 3'b110;
        rom_memory[45982] = 3'b110;
        rom_memory[45983] = 3'b110;
        rom_memory[45984] = 3'b110;
        rom_memory[45985] = 3'b110;
        rom_memory[45986] = 3'b110;
        rom_memory[45987] = 3'b110;
        rom_memory[45988] = 3'b110;
        rom_memory[45989] = 3'b110;
        rom_memory[45990] = 3'b110;
        rom_memory[45991] = 3'b110;
        rom_memory[45992] = 3'b110;
        rom_memory[45993] = 3'b110;
        rom_memory[45994] = 3'b110;
        rom_memory[45995] = 3'b110;
        rom_memory[45996] = 3'b110;
        rom_memory[45997] = 3'b110;
        rom_memory[45998] = 3'b110;
        rom_memory[45999] = 3'b110;
        rom_memory[46000] = 3'b110;
        rom_memory[46001] = 3'b110;
        rom_memory[46002] = 3'b110;
        rom_memory[46003] = 3'b110;
        rom_memory[46004] = 3'b110;
        rom_memory[46005] = 3'b110;
        rom_memory[46006] = 3'b110;
        rom_memory[46007] = 3'b110;
        rom_memory[46008] = 3'b110;
        rom_memory[46009] = 3'b110;
        rom_memory[46010] = 3'b110;
        rom_memory[46011] = 3'b110;
        rom_memory[46012] = 3'b110;
        rom_memory[46013] = 3'b110;
        rom_memory[46014] = 3'b110;
        rom_memory[46015] = 3'b110;
        rom_memory[46016] = 3'b110;
        rom_memory[46017] = 3'b110;
        rom_memory[46018] = 3'b110;
        rom_memory[46019] = 3'b110;
        rom_memory[46020] = 3'b110;
        rom_memory[46021] = 3'b110;
        rom_memory[46022] = 3'b110;
        rom_memory[46023] = 3'b110;
        rom_memory[46024] = 3'b110;
        rom_memory[46025] = 3'b110;
        rom_memory[46026] = 3'b110;
        rom_memory[46027] = 3'b110;
        rom_memory[46028] = 3'b110;
        rom_memory[46029] = 3'b110;
        rom_memory[46030] = 3'b110;
        rom_memory[46031] = 3'b110;
        rom_memory[46032] = 3'b110;
        rom_memory[46033] = 3'b110;
        rom_memory[46034] = 3'b110;
        rom_memory[46035] = 3'b110;
        rom_memory[46036] = 3'b110;
        rom_memory[46037] = 3'b110;
        rom_memory[46038] = 3'b110;
        rom_memory[46039] = 3'b110;
        rom_memory[46040] = 3'b110;
        rom_memory[46041] = 3'b110;
        rom_memory[46042] = 3'b110;
        rom_memory[46043] = 3'b110;
        rom_memory[46044] = 3'b110;
        rom_memory[46045] = 3'b110;
        rom_memory[46046] = 3'b110;
        rom_memory[46047] = 3'b110;
        rom_memory[46048] = 3'b110;
        rom_memory[46049] = 3'b110;
        rom_memory[46050] = 3'b100;
        rom_memory[46051] = 3'b000;
        rom_memory[46052] = 3'b000;
        rom_memory[46053] = 3'b000;
        rom_memory[46054] = 3'b000;
        rom_memory[46055] = 3'b000;
        rom_memory[46056] = 3'b000;
        rom_memory[46057] = 3'b000;
        rom_memory[46058] = 3'b110;
        rom_memory[46059] = 3'b110;
        rom_memory[46060] = 3'b110;
        rom_memory[46061] = 3'b110;
        rom_memory[46062] = 3'b110;
        rom_memory[46063] = 3'b110;
        rom_memory[46064] = 3'b110;
        rom_memory[46065] = 3'b110;
        rom_memory[46066] = 3'b110;
        rom_memory[46067] = 3'b110;
        rom_memory[46068] = 3'b110;
        rom_memory[46069] = 3'b110;
        rom_memory[46070] = 3'b110;
        rom_memory[46071] = 3'b110;
        rom_memory[46072] = 3'b110;
        rom_memory[46073] = 3'b110;
        rom_memory[46074] = 3'b110;
        rom_memory[46075] = 3'b110;
        rom_memory[46076] = 3'b110;
        rom_memory[46077] = 3'b110;
        rom_memory[46078] = 3'b110;
        rom_memory[46079] = 3'b110;
        rom_memory[46080] = 3'b111;
        rom_memory[46081] = 3'b111;
        rom_memory[46082] = 3'b111;
        rom_memory[46083] = 3'b111;
        rom_memory[46084] = 3'b111;
        rom_memory[46085] = 3'b111;
        rom_memory[46086] = 3'b111;
        rom_memory[46087] = 3'b111;
        rom_memory[46088] = 3'b111;
        rom_memory[46089] = 3'b111;
        rom_memory[46090] = 3'b111;
        rom_memory[46091] = 3'b111;
        rom_memory[46092] = 3'b111;
        rom_memory[46093] = 3'b111;
        rom_memory[46094] = 3'b111;
        rom_memory[46095] = 3'b111;
        rom_memory[46096] = 3'b111;
        rom_memory[46097] = 3'b111;
        rom_memory[46098] = 3'b111;
        rom_memory[46099] = 3'b111;
        rom_memory[46100] = 3'b110;
        rom_memory[46101] = 3'b110;
        rom_memory[46102] = 3'b110;
        rom_memory[46103] = 3'b110;
        rom_memory[46104] = 3'b110;
        rom_memory[46105] = 3'b110;
        rom_memory[46106] = 3'b110;
        rom_memory[46107] = 3'b110;
        rom_memory[46108] = 3'b110;
        rom_memory[46109] = 3'b110;
        rom_memory[46110] = 3'b111;
        rom_memory[46111] = 3'b111;
        rom_memory[46112] = 3'b111;
        rom_memory[46113] = 3'b111;
        rom_memory[46114] = 3'b111;
        rom_memory[46115] = 3'b111;
        rom_memory[46116] = 3'b111;
        rom_memory[46117] = 3'b111;
        rom_memory[46118] = 3'b111;
        rom_memory[46119] = 3'b111;
        rom_memory[46120] = 3'b111;
        rom_memory[46121] = 3'b111;
        rom_memory[46122] = 3'b111;
        rom_memory[46123] = 3'b111;
        rom_memory[46124] = 3'b111;
        rom_memory[46125] = 3'b111;
        rom_memory[46126] = 3'b111;
        rom_memory[46127] = 3'b111;
        rom_memory[46128] = 3'b111;
        rom_memory[46129] = 3'b111;
        rom_memory[46130] = 3'b110;
        rom_memory[46131] = 3'b110;
        rom_memory[46132] = 3'b110;
        rom_memory[46133] = 3'b110;
        rom_memory[46134] = 3'b111;
        rom_memory[46135] = 3'b111;
        rom_memory[46136] = 3'b110;
        rom_memory[46137] = 3'b110;
        rom_memory[46138] = 3'b100;
        rom_memory[46139] = 3'b100;
        rom_memory[46140] = 3'b100;
        rom_memory[46141] = 3'b000;
        rom_memory[46142] = 3'b000;
        rom_memory[46143] = 3'b100;
        rom_memory[46144] = 3'b110;
        rom_memory[46145] = 3'b111;
        rom_memory[46146] = 3'b111;
        rom_memory[46147] = 3'b111;
        rom_memory[46148] = 3'b111;
        rom_memory[46149] = 3'b111;
        rom_memory[46150] = 3'b111;
        rom_memory[46151] = 3'b100;
        rom_memory[46152] = 3'b110;
        rom_memory[46153] = 3'b000;
        rom_memory[46154] = 3'b000;
        rom_memory[46155] = 3'b111;
        rom_memory[46156] = 3'b111;
        rom_memory[46157] = 3'b111;
        rom_memory[46158] = 3'b110;
        rom_memory[46159] = 3'b111;
        rom_memory[46160] = 3'b110;
        rom_memory[46161] = 3'b110;
        rom_memory[46162] = 3'b111;
        rom_memory[46163] = 3'b111;
        rom_memory[46164] = 3'b111;
        rom_memory[46165] = 3'b111;
        rom_memory[46166] = 3'b111;
        rom_memory[46167] = 3'b111;
        rom_memory[46168] = 3'b100;
        rom_memory[46169] = 3'b110;
        rom_memory[46170] = 3'b100;
        rom_memory[46171] = 3'b110;
        rom_memory[46172] = 3'b111;
        rom_memory[46173] = 3'b111;
        rom_memory[46174] = 3'b110;
        rom_memory[46175] = 3'b110;
        rom_memory[46176] = 3'b110;
        rom_memory[46177] = 3'b110;
        rom_memory[46178] = 3'b110;
        rom_memory[46179] = 3'b110;
        rom_memory[46180] = 3'b110;
        rom_memory[46181] = 3'b110;
        rom_memory[46182] = 3'b110;
        rom_memory[46183] = 3'b110;
        rom_memory[46184] = 3'b111;
        rom_memory[46185] = 3'b111;
        rom_memory[46186] = 3'b111;
        rom_memory[46187] = 3'b111;
        rom_memory[46188] = 3'b111;
        rom_memory[46189] = 3'b111;
        rom_memory[46190] = 3'b111;
        rom_memory[46191] = 3'b111;
        rom_memory[46192] = 3'b111;
        rom_memory[46193] = 3'b111;
        rom_memory[46194] = 3'b111;
        rom_memory[46195] = 3'b111;
        rom_memory[46196] = 3'b111;
        rom_memory[46197] = 3'b110;
        rom_memory[46198] = 3'b110;
        rom_memory[46199] = 3'b110;
        rom_memory[46200] = 3'b110;
        rom_memory[46201] = 3'b110;
        rom_memory[46202] = 3'b110;
        rom_memory[46203] = 3'b110;
        rom_memory[46204] = 3'b110;
        rom_memory[46205] = 3'b110;
        rom_memory[46206] = 3'b110;
        rom_memory[46207] = 3'b110;
        rom_memory[46208] = 3'b110;
        rom_memory[46209] = 3'b110;
        rom_memory[46210] = 3'b110;
        rom_memory[46211] = 3'b110;
        rom_memory[46212] = 3'b110;
        rom_memory[46213] = 3'b110;
        rom_memory[46214] = 3'b110;
        rom_memory[46215] = 3'b110;
        rom_memory[46216] = 3'b110;
        rom_memory[46217] = 3'b110;
        rom_memory[46218] = 3'b110;
        rom_memory[46219] = 3'b110;
        rom_memory[46220] = 3'b110;
        rom_memory[46221] = 3'b110;
        rom_memory[46222] = 3'b110;
        rom_memory[46223] = 3'b110;
        rom_memory[46224] = 3'b110;
        rom_memory[46225] = 3'b110;
        rom_memory[46226] = 3'b110;
        rom_memory[46227] = 3'b110;
        rom_memory[46228] = 3'b110;
        rom_memory[46229] = 3'b110;
        rom_memory[46230] = 3'b110;
        rom_memory[46231] = 3'b110;
        rom_memory[46232] = 3'b110;
        rom_memory[46233] = 3'b110;
        rom_memory[46234] = 3'b110;
        rom_memory[46235] = 3'b110;
        rom_memory[46236] = 3'b110;
        rom_memory[46237] = 3'b110;
        rom_memory[46238] = 3'b110;
        rom_memory[46239] = 3'b110;
        rom_memory[46240] = 3'b110;
        rom_memory[46241] = 3'b110;
        rom_memory[46242] = 3'b110;
        rom_memory[46243] = 3'b110;
        rom_memory[46244] = 3'b110;
        rom_memory[46245] = 3'b110;
        rom_memory[46246] = 3'b110;
        rom_memory[46247] = 3'b110;
        rom_memory[46248] = 3'b110;
        rom_memory[46249] = 3'b110;
        rom_memory[46250] = 3'b110;
        rom_memory[46251] = 3'b110;
        rom_memory[46252] = 3'b110;
        rom_memory[46253] = 3'b110;
        rom_memory[46254] = 3'b110;
        rom_memory[46255] = 3'b110;
        rom_memory[46256] = 3'b110;
        rom_memory[46257] = 3'b110;
        rom_memory[46258] = 3'b110;
        rom_memory[46259] = 3'b110;
        rom_memory[46260] = 3'b110;
        rom_memory[46261] = 3'b110;
        rom_memory[46262] = 3'b110;
        rom_memory[46263] = 3'b110;
        rom_memory[46264] = 3'b110;
        rom_memory[46265] = 3'b110;
        rom_memory[46266] = 3'b110;
        rom_memory[46267] = 3'b110;
        rom_memory[46268] = 3'b110;
        rom_memory[46269] = 3'b110;
        rom_memory[46270] = 3'b110;
        rom_memory[46271] = 3'b110;
        rom_memory[46272] = 3'b110;
        rom_memory[46273] = 3'b110;
        rom_memory[46274] = 3'b110;
        rom_memory[46275] = 3'b110;
        rom_memory[46276] = 3'b110;
        rom_memory[46277] = 3'b110;
        rom_memory[46278] = 3'b110;
        rom_memory[46279] = 3'b110;
        rom_memory[46280] = 3'b110;
        rom_memory[46281] = 3'b110;
        rom_memory[46282] = 3'b110;
        rom_memory[46283] = 3'b110;
        rom_memory[46284] = 3'b110;
        rom_memory[46285] = 3'b110;
        rom_memory[46286] = 3'b110;
        rom_memory[46287] = 3'b110;
        rom_memory[46288] = 3'b110;
        rom_memory[46289] = 3'b110;
        rom_memory[46290] = 3'b110;
        rom_memory[46291] = 3'b110;
        rom_memory[46292] = 3'b000;
        rom_memory[46293] = 3'b000;
        rom_memory[46294] = 3'b000;
        rom_memory[46295] = 3'b000;
        rom_memory[46296] = 3'b000;
        rom_memory[46297] = 3'b000;
        rom_memory[46298] = 3'b000;
        rom_memory[46299] = 3'b100;
        rom_memory[46300] = 3'b110;
        rom_memory[46301] = 3'b110;
        rom_memory[46302] = 3'b110;
        rom_memory[46303] = 3'b110;
        rom_memory[46304] = 3'b110;
        rom_memory[46305] = 3'b110;
        rom_memory[46306] = 3'b110;
        rom_memory[46307] = 3'b110;
        rom_memory[46308] = 3'b110;
        rom_memory[46309] = 3'b110;
        rom_memory[46310] = 3'b110;
        rom_memory[46311] = 3'b110;
        rom_memory[46312] = 3'b110;
        rom_memory[46313] = 3'b110;
        rom_memory[46314] = 3'b110;
        rom_memory[46315] = 3'b110;
        rom_memory[46316] = 3'b110;
        rom_memory[46317] = 3'b110;
        rom_memory[46318] = 3'b110;
        rom_memory[46319] = 3'b110;
        rom_memory[46320] = 3'b111;
        rom_memory[46321] = 3'b111;
        rom_memory[46322] = 3'b111;
        rom_memory[46323] = 3'b111;
        rom_memory[46324] = 3'b111;
        rom_memory[46325] = 3'b111;
        rom_memory[46326] = 3'b111;
        rom_memory[46327] = 3'b111;
        rom_memory[46328] = 3'b111;
        rom_memory[46329] = 3'b111;
        rom_memory[46330] = 3'b111;
        rom_memory[46331] = 3'b111;
        rom_memory[46332] = 3'b111;
        rom_memory[46333] = 3'b111;
        rom_memory[46334] = 3'b111;
        rom_memory[46335] = 3'b111;
        rom_memory[46336] = 3'b111;
        rom_memory[46337] = 3'b111;
        rom_memory[46338] = 3'b111;
        rom_memory[46339] = 3'b110;
        rom_memory[46340] = 3'b110;
        rom_memory[46341] = 3'b110;
        rom_memory[46342] = 3'b110;
        rom_memory[46343] = 3'b110;
        rom_memory[46344] = 3'b110;
        rom_memory[46345] = 3'b110;
        rom_memory[46346] = 3'b110;
        rom_memory[46347] = 3'b110;
        rom_memory[46348] = 3'b110;
        rom_memory[46349] = 3'b110;
        rom_memory[46350] = 3'b110;
        rom_memory[46351] = 3'b111;
        rom_memory[46352] = 3'b111;
        rom_memory[46353] = 3'b111;
        rom_memory[46354] = 3'b111;
        rom_memory[46355] = 3'b111;
        rom_memory[46356] = 3'b111;
        rom_memory[46357] = 3'b111;
        rom_memory[46358] = 3'b111;
        rom_memory[46359] = 3'b111;
        rom_memory[46360] = 3'b111;
        rom_memory[46361] = 3'b111;
        rom_memory[46362] = 3'b111;
        rom_memory[46363] = 3'b110;
        rom_memory[46364] = 3'b111;
        rom_memory[46365] = 3'b111;
        rom_memory[46366] = 3'b111;
        rom_memory[46367] = 3'b111;
        rom_memory[46368] = 3'b111;
        rom_memory[46369] = 3'b111;
        rom_memory[46370] = 3'b110;
        rom_memory[46371] = 3'b110;
        rom_memory[46372] = 3'b110;
        rom_memory[46373] = 3'b110;
        rom_memory[46374] = 3'b111;
        rom_memory[46375] = 3'b111;
        rom_memory[46376] = 3'b110;
        rom_memory[46377] = 3'b110;
        rom_memory[46378] = 3'b100;
        rom_memory[46379] = 3'b100;
        rom_memory[46380] = 3'b000;
        rom_memory[46381] = 3'b000;
        rom_memory[46382] = 3'b000;
        rom_memory[46383] = 3'b100;
        rom_memory[46384] = 3'b100;
        rom_memory[46385] = 3'b111;
        rom_memory[46386] = 3'b111;
        rom_memory[46387] = 3'b111;
        rom_memory[46388] = 3'b111;
        rom_memory[46389] = 3'b111;
        rom_memory[46390] = 3'b111;
        rom_memory[46391] = 3'b110;
        rom_memory[46392] = 3'b100;
        rom_memory[46393] = 3'b000;
        rom_memory[46394] = 3'b000;
        rom_memory[46395] = 3'b111;
        rom_memory[46396] = 3'b111;
        rom_memory[46397] = 3'b111;
        rom_memory[46398] = 3'b111;
        rom_memory[46399] = 3'b111;
        rom_memory[46400] = 3'b100;
        rom_memory[46401] = 3'b100;
        rom_memory[46402] = 3'b111;
        rom_memory[46403] = 3'b110;
        rom_memory[46404] = 3'b110;
        rom_memory[46405] = 3'b100;
        rom_memory[46406] = 3'b000;
        rom_memory[46407] = 3'b000;
        rom_memory[46408] = 3'b100;
        rom_memory[46409] = 3'b111;
        rom_memory[46410] = 3'b100;
        rom_memory[46411] = 3'b111;
        rom_memory[46412] = 3'b111;
        rom_memory[46413] = 3'b111;
        rom_memory[46414] = 3'b111;
        rom_memory[46415] = 3'b110;
        rom_memory[46416] = 3'b110;
        rom_memory[46417] = 3'b110;
        rom_memory[46418] = 3'b110;
        rom_memory[46419] = 3'b110;
        rom_memory[46420] = 3'b110;
        rom_memory[46421] = 3'b110;
        rom_memory[46422] = 3'b110;
        rom_memory[46423] = 3'b111;
        rom_memory[46424] = 3'b111;
        rom_memory[46425] = 3'b111;
        rom_memory[46426] = 3'b111;
        rom_memory[46427] = 3'b111;
        rom_memory[46428] = 3'b111;
        rom_memory[46429] = 3'b111;
        rom_memory[46430] = 3'b111;
        rom_memory[46431] = 3'b111;
        rom_memory[46432] = 3'b111;
        rom_memory[46433] = 3'b111;
        rom_memory[46434] = 3'b111;
        rom_memory[46435] = 3'b111;
        rom_memory[46436] = 3'b111;
        rom_memory[46437] = 3'b110;
        rom_memory[46438] = 3'b110;
        rom_memory[46439] = 3'b110;
        rom_memory[46440] = 3'b110;
        rom_memory[46441] = 3'b110;
        rom_memory[46442] = 3'b110;
        rom_memory[46443] = 3'b110;
        rom_memory[46444] = 3'b110;
        rom_memory[46445] = 3'b110;
        rom_memory[46446] = 3'b110;
        rom_memory[46447] = 3'b110;
        rom_memory[46448] = 3'b110;
        rom_memory[46449] = 3'b110;
        rom_memory[46450] = 3'b110;
        rom_memory[46451] = 3'b110;
        rom_memory[46452] = 3'b110;
        rom_memory[46453] = 3'b110;
        rom_memory[46454] = 3'b110;
        rom_memory[46455] = 3'b110;
        rom_memory[46456] = 3'b110;
        rom_memory[46457] = 3'b110;
        rom_memory[46458] = 3'b110;
        rom_memory[46459] = 3'b110;
        rom_memory[46460] = 3'b110;
        rom_memory[46461] = 3'b110;
        rom_memory[46462] = 3'b110;
        rom_memory[46463] = 3'b110;
        rom_memory[46464] = 3'b110;
        rom_memory[46465] = 3'b110;
        rom_memory[46466] = 3'b110;
        rom_memory[46467] = 3'b110;
        rom_memory[46468] = 3'b110;
        rom_memory[46469] = 3'b110;
        rom_memory[46470] = 3'b110;
        rom_memory[46471] = 3'b110;
        rom_memory[46472] = 3'b110;
        rom_memory[46473] = 3'b110;
        rom_memory[46474] = 3'b110;
        rom_memory[46475] = 3'b110;
        rom_memory[46476] = 3'b110;
        rom_memory[46477] = 3'b110;
        rom_memory[46478] = 3'b110;
        rom_memory[46479] = 3'b110;
        rom_memory[46480] = 3'b110;
        rom_memory[46481] = 3'b110;
        rom_memory[46482] = 3'b110;
        rom_memory[46483] = 3'b110;
        rom_memory[46484] = 3'b110;
        rom_memory[46485] = 3'b110;
        rom_memory[46486] = 3'b110;
        rom_memory[46487] = 3'b110;
        rom_memory[46488] = 3'b110;
        rom_memory[46489] = 3'b110;
        rom_memory[46490] = 3'b110;
        rom_memory[46491] = 3'b110;
        rom_memory[46492] = 3'b110;
        rom_memory[46493] = 3'b110;
        rom_memory[46494] = 3'b110;
        rom_memory[46495] = 3'b110;
        rom_memory[46496] = 3'b110;
        rom_memory[46497] = 3'b110;
        rom_memory[46498] = 3'b110;
        rom_memory[46499] = 3'b110;
        rom_memory[46500] = 3'b110;
        rom_memory[46501] = 3'b110;
        rom_memory[46502] = 3'b110;
        rom_memory[46503] = 3'b110;
        rom_memory[46504] = 3'b110;
        rom_memory[46505] = 3'b110;
        rom_memory[46506] = 3'b110;
        rom_memory[46507] = 3'b110;
        rom_memory[46508] = 3'b110;
        rom_memory[46509] = 3'b110;
        rom_memory[46510] = 3'b110;
        rom_memory[46511] = 3'b110;
        rom_memory[46512] = 3'b110;
        rom_memory[46513] = 3'b110;
        rom_memory[46514] = 3'b110;
        rom_memory[46515] = 3'b110;
        rom_memory[46516] = 3'b110;
        rom_memory[46517] = 3'b110;
        rom_memory[46518] = 3'b110;
        rom_memory[46519] = 3'b110;
        rom_memory[46520] = 3'b110;
        rom_memory[46521] = 3'b110;
        rom_memory[46522] = 3'b110;
        rom_memory[46523] = 3'b110;
        rom_memory[46524] = 3'b110;
        rom_memory[46525] = 3'b110;
        rom_memory[46526] = 3'b110;
        rom_memory[46527] = 3'b110;
        rom_memory[46528] = 3'b110;
        rom_memory[46529] = 3'b110;
        rom_memory[46530] = 3'b110;
        rom_memory[46531] = 3'b110;
        rom_memory[46532] = 3'b110;
        rom_memory[46533] = 3'b110;
        rom_memory[46534] = 3'b100;
        rom_memory[46535] = 3'b000;
        rom_memory[46536] = 3'b000;
        rom_memory[46537] = 3'b000;
        rom_memory[46538] = 3'b000;
        rom_memory[46539] = 3'b000;
        rom_memory[46540] = 3'b000;
        rom_memory[46541] = 3'b110;
        rom_memory[46542] = 3'b110;
        rom_memory[46543] = 3'b110;
        rom_memory[46544] = 3'b110;
        rom_memory[46545] = 3'b110;
        rom_memory[46546] = 3'b110;
        rom_memory[46547] = 3'b110;
        rom_memory[46548] = 3'b110;
        rom_memory[46549] = 3'b110;
        rom_memory[46550] = 3'b110;
        rom_memory[46551] = 3'b110;
        rom_memory[46552] = 3'b110;
        rom_memory[46553] = 3'b110;
        rom_memory[46554] = 3'b110;
        rom_memory[46555] = 3'b110;
        rom_memory[46556] = 3'b110;
        rom_memory[46557] = 3'b110;
        rom_memory[46558] = 3'b110;
        rom_memory[46559] = 3'b110;
        rom_memory[46560] = 3'b111;
        rom_memory[46561] = 3'b111;
        rom_memory[46562] = 3'b111;
        rom_memory[46563] = 3'b111;
        rom_memory[46564] = 3'b111;
        rom_memory[46565] = 3'b111;
        rom_memory[46566] = 3'b111;
        rom_memory[46567] = 3'b111;
        rom_memory[46568] = 3'b111;
        rom_memory[46569] = 3'b111;
        rom_memory[46570] = 3'b111;
        rom_memory[46571] = 3'b111;
        rom_memory[46572] = 3'b111;
        rom_memory[46573] = 3'b111;
        rom_memory[46574] = 3'b111;
        rom_memory[46575] = 3'b111;
        rom_memory[46576] = 3'b111;
        rom_memory[46577] = 3'b111;
        rom_memory[46578] = 3'b111;
        rom_memory[46579] = 3'b110;
        rom_memory[46580] = 3'b110;
        rom_memory[46581] = 3'b110;
        rom_memory[46582] = 3'b110;
        rom_memory[46583] = 3'b110;
        rom_memory[46584] = 3'b110;
        rom_memory[46585] = 3'b110;
        rom_memory[46586] = 3'b110;
        rom_memory[46587] = 3'b110;
        rom_memory[46588] = 3'b110;
        rom_memory[46589] = 3'b110;
        rom_memory[46590] = 3'b110;
        rom_memory[46591] = 3'b111;
        rom_memory[46592] = 3'b111;
        rom_memory[46593] = 3'b111;
        rom_memory[46594] = 3'b111;
        rom_memory[46595] = 3'b111;
        rom_memory[46596] = 3'b111;
        rom_memory[46597] = 3'b111;
        rom_memory[46598] = 3'b111;
        rom_memory[46599] = 3'b110;
        rom_memory[46600] = 3'b110;
        rom_memory[46601] = 3'b110;
        rom_memory[46602] = 3'b111;
        rom_memory[46603] = 3'b111;
        rom_memory[46604] = 3'b110;
        rom_memory[46605] = 3'b111;
        rom_memory[46606] = 3'b111;
        rom_memory[46607] = 3'b111;
        rom_memory[46608] = 3'b111;
        rom_memory[46609] = 3'b111;
        rom_memory[46610] = 3'b110;
        rom_memory[46611] = 3'b110;
        rom_memory[46612] = 3'b110;
        rom_memory[46613] = 3'b110;
        rom_memory[46614] = 3'b111;
        rom_memory[46615] = 3'b110;
        rom_memory[46616] = 3'b110;
        rom_memory[46617] = 3'b110;
        rom_memory[46618] = 3'b110;
        rom_memory[46619] = 3'b100;
        rom_memory[46620] = 3'b100;
        rom_memory[46621] = 3'b000;
        rom_memory[46622] = 3'b000;
        rom_memory[46623] = 3'b100;
        rom_memory[46624] = 3'b000;
        rom_memory[46625] = 3'b111;
        rom_memory[46626] = 3'b100;
        rom_memory[46627] = 3'b110;
        rom_memory[46628] = 3'b110;
        rom_memory[46629] = 3'b111;
        rom_memory[46630] = 3'b111;
        rom_memory[46631] = 3'b110;
        rom_memory[46632] = 3'b100;
        rom_memory[46633] = 3'b000;
        rom_memory[46634] = 3'b000;
        rom_memory[46635] = 3'b111;
        rom_memory[46636] = 3'b000;
        rom_memory[46637] = 3'b100;
        rom_memory[46638] = 3'b111;
        rom_memory[46639] = 3'b000;
        rom_memory[46640] = 3'b111;
        rom_memory[46641] = 3'b111;
        rom_memory[46642] = 3'b000;
        rom_memory[46643] = 3'b111;
        rom_memory[46644] = 3'b110;
        rom_memory[46645] = 3'b000;
        rom_memory[46646] = 3'b000;
        rom_memory[46647] = 3'b000;
        rom_memory[46648] = 3'b000;
        rom_memory[46649] = 3'b111;
        rom_memory[46650] = 3'b111;
        rom_memory[46651] = 3'b111;
        rom_memory[46652] = 3'b111;
        rom_memory[46653] = 3'b111;
        rom_memory[46654] = 3'b111;
        rom_memory[46655] = 3'b110;
        rom_memory[46656] = 3'b110;
        rom_memory[46657] = 3'b110;
        rom_memory[46658] = 3'b110;
        rom_memory[46659] = 3'b110;
        rom_memory[46660] = 3'b110;
        rom_memory[46661] = 3'b110;
        rom_memory[46662] = 3'b110;
        rom_memory[46663] = 3'b111;
        rom_memory[46664] = 3'b111;
        rom_memory[46665] = 3'b111;
        rom_memory[46666] = 3'b111;
        rom_memory[46667] = 3'b111;
        rom_memory[46668] = 3'b111;
        rom_memory[46669] = 3'b111;
        rom_memory[46670] = 3'b111;
        rom_memory[46671] = 3'b111;
        rom_memory[46672] = 3'b111;
        rom_memory[46673] = 3'b111;
        rom_memory[46674] = 3'b111;
        rom_memory[46675] = 3'b111;
        rom_memory[46676] = 3'b111;
        rom_memory[46677] = 3'b110;
        rom_memory[46678] = 3'b110;
        rom_memory[46679] = 3'b110;
        rom_memory[46680] = 3'b110;
        rom_memory[46681] = 3'b110;
        rom_memory[46682] = 3'b110;
        rom_memory[46683] = 3'b110;
        rom_memory[46684] = 3'b110;
        rom_memory[46685] = 3'b110;
        rom_memory[46686] = 3'b110;
        rom_memory[46687] = 3'b110;
        rom_memory[46688] = 3'b110;
        rom_memory[46689] = 3'b110;
        rom_memory[46690] = 3'b110;
        rom_memory[46691] = 3'b110;
        rom_memory[46692] = 3'b110;
        rom_memory[46693] = 3'b110;
        rom_memory[46694] = 3'b110;
        rom_memory[46695] = 3'b110;
        rom_memory[46696] = 3'b110;
        rom_memory[46697] = 3'b110;
        rom_memory[46698] = 3'b110;
        rom_memory[46699] = 3'b110;
        rom_memory[46700] = 3'b110;
        rom_memory[46701] = 3'b110;
        rom_memory[46702] = 3'b110;
        rom_memory[46703] = 3'b110;
        rom_memory[46704] = 3'b110;
        rom_memory[46705] = 3'b110;
        rom_memory[46706] = 3'b110;
        rom_memory[46707] = 3'b110;
        rom_memory[46708] = 3'b110;
        rom_memory[46709] = 3'b110;
        rom_memory[46710] = 3'b110;
        rom_memory[46711] = 3'b110;
        rom_memory[46712] = 3'b110;
        rom_memory[46713] = 3'b110;
        rom_memory[46714] = 3'b110;
        rom_memory[46715] = 3'b110;
        rom_memory[46716] = 3'b110;
        rom_memory[46717] = 3'b110;
        rom_memory[46718] = 3'b110;
        rom_memory[46719] = 3'b110;
        rom_memory[46720] = 3'b110;
        rom_memory[46721] = 3'b110;
        rom_memory[46722] = 3'b110;
        rom_memory[46723] = 3'b110;
        rom_memory[46724] = 3'b110;
        rom_memory[46725] = 3'b110;
        rom_memory[46726] = 3'b110;
        rom_memory[46727] = 3'b110;
        rom_memory[46728] = 3'b110;
        rom_memory[46729] = 3'b110;
        rom_memory[46730] = 3'b110;
        rom_memory[46731] = 3'b110;
        rom_memory[46732] = 3'b110;
        rom_memory[46733] = 3'b110;
        rom_memory[46734] = 3'b110;
        rom_memory[46735] = 3'b110;
        rom_memory[46736] = 3'b110;
        rom_memory[46737] = 3'b110;
        rom_memory[46738] = 3'b110;
        rom_memory[46739] = 3'b110;
        rom_memory[46740] = 3'b110;
        rom_memory[46741] = 3'b110;
        rom_memory[46742] = 3'b110;
        rom_memory[46743] = 3'b110;
        rom_memory[46744] = 3'b110;
        rom_memory[46745] = 3'b110;
        rom_memory[46746] = 3'b110;
        rom_memory[46747] = 3'b110;
        rom_memory[46748] = 3'b110;
        rom_memory[46749] = 3'b110;
        rom_memory[46750] = 3'b110;
        rom_memory[46751] = 3'b110;
        rom_memory[46752] = 3'b110;
        rom_memory[46753] = 3'b110;
        rom_memory[46754] = 3'b110;
        rom_memory[46755] = 3'b110;
        rom_memory[46756] = 3'b110;
        rom_memory[46757] = 3'b110;
        rom_memory[46758] = 3'b110;
        rom_memory[46759] = 3'b110;
        rom_memory[46760] = 3'b110;
        rom_memory[46761] = 3'b110;
        rom_memory[46762] = 3'b110;
        rom_memory[46763] = 3'b110;
        rom_memory[46764] = 3'b110;
        rom_memory[46765] = 3'b110;
        rom_memory[46766] = 3'b110;
        rom_memory[46767] = 3'b110;
        rom_memory[46768] = 3'b110;
        rom_memory[46769] = 3'b110;
        rom_memory[46770] = 3'b110;
        rom_memory[46771] = 3'b110;
        rom_memory[46772] = 3'b110;
        rom_memory[46773] = 3'b110;
        rom_memory[46774] = 3'b110;
        rom_memory[46775] = 3'b110;
        rom_memory[46776] = 3'b100;
        rom_memory[46777] = 3'b000;
        rom_memory[46778] = 3'b000;
        rom_memory[46779] = 3'b000;
        rom_memory[46780] = 3'b000;
        rom_memory[46781] = 3'b000;
        rom_memory[46782] = 3'b000;
        rom_memory[46783] = 3'b110;
        rom_memory[46784] = 3'b110;
        rom_memory[46785] = 3'b110;
        rom_memory[46786] = 3'b110;
        rom_memory[46787] = 3'b110;
        rom_memory[46788] = 3'b110;
        rom_memory[46789] = 3'b110;
        rom_memory[46790] = 3'b110;
        rom_memory[46791] = 3'b110;
        rom_memory[46792] = 3'b110;
        rom_memory[46793] = 3'b110;
        rom_memory[46794] = 3'b110;
        rom_memory[46795] = 3'b110;
        rom_memory[46796] = 3'b110;
        rom_memory[46797] = 3'b110;
        rom_memory[46798] = 3'b110;
        rom_memory[46799] = 3'b110;
        rom_memory[46800] = 3'b111;
        rom_memory[46801] = 3'b111;
        rom_memory[46802] = 3'b111;
        rom_memory[46803] = 3'b111;
        rom_memory[46804] = 3'b111;
        rom_memory[46805] = 3'b111;
        rom_memory[46806] = 3'b111;
        rom_memory[46807] = 3'b111;
        rom_memory[46808] = 3'b111;
        rom_memory[46809] = 3'b111;
        rom_memory[46810] = 3'b111;
        rom_memory[46811] = 3'b111;
        rom_memory[46812] = 3'b111;
        rom_memory[46813] = 3'b111;
        rom_memory[46814] = 3'b111;
        rom_memory[46815] = 3'b111;
        rom_memory[46816] = 3'b111;
        rom_memory[46817] = 3'b111;
        rom_memory[46818] = 3'b110;
        rom_memory[46819] = 3'b110;
        rom_memory[46820] = 3'b110;
        rom_memory[46821] = 3'b110;
        rom_memory[46822] = 3'b110;
        rom_memory[46823] = 3'b110;
        rom_memory[46824] = 3'b110;
        rom_memory[46825] = 3'b110;
        rom_memory[46826] = 3'b110;
        rom_memory[46827] = 3'b110;
        rom_memory[46828] = 3'b110;
        rom_memory[46829] = 3'b110;
        rom_memory[46830] = 3'b110;
        rom_memory[46831] = 3'b111;
        rom_memory[46832] = 3'b111;
        rom_memory[46833] = 3'b111;
        rom_memory[46834] = 3'b111;
        rom_memory[46835] = 3'b111;
        rom_memory[46836] = 3'b111;
        rom_memory[46837] = 3'b111;
        rom_memory[46838] = 3'b110;
        rom_memory[46839] = 3'b110;
        rom_memory[46840] = 3'b110;
        rom_memory[46841] = 3'b110;
        rom_memory[46842] = 3'b111;
        rom_memory[46843] = 3'b111;
        rom_memory[46844] = 3'b111;
        rom_memory[46845] = 3'b110;
        rom_memory[46846] = 3'b111;
        rom_memory[46847] = 3'b111;
        rom_memory[46848] = 3'b111;
        rom_memory[46849] = 3'b111;
        rom_memory[46850] = 3'b110;
        rom_memory[46851] = 3'b110;
        rom_memory[46852] = 3'b110;
        rom_memory[46853] = 3'b110;
        rom_memory[46854] = 3'b110;
        rom_memory[46855] = 3'b110;
        rom_memory[46856] = 3'b110;
        rom_memory[46857] = 3'b110;
        rom_memory[46858] = 3'b110;
        rom_memory[46859] = 3'b110;
        rom_memory[46860] = 3'b100;
        rom_memory[46861] = 3'b100;
        rom_memory[46862] = 3'b100;
        rom_memory[46863] = 3'b110;
        rom_memory[46864] = 3'b100;
        rom_memory[46865] = 3'b100;
        rom_memory[46866] = 3'b111;
        rom_memory[46867] = 3'b111;
        rom_memory[46868] = 3'b110;
        rom_memory[46869] = 3'b111;
        rom_memory[46870] = 3'b111;
        rom_memory[46871] = 3'b110;
        rom_memory[46872] = 3'b111;
        rom_memory[46873] = 3'b000;
        rom_memory[46874] = 3'b000;
        rom_memory[46875] = 3'b100;
        rom_memory[46876] = 3'b000;
        rom_memory[46877] = 3'b000;
        rom_memory[46878] = 3'b100;
        rom_memory[46879] = 3'b100;
        rom_memory[46880] = 3'b000;
        rom_memory[46881] = 3'b110;
        rom_memory[46882] = 3'b100;
        rom_memory[46883] = 3'b000;
        rom_memory[46884] = 3'b100;
        rom_memory[46885] = 3'b100;
        rom_memory[46886] = 3'b100;
        rom_memory[46887] = 3'b111;
        rom_memory[46888] = 3'b110;
        rom_memory[46889] = 3'b100;
        rom_memory[46890] = 3'b111;
        rom_memory[46891] = 3'b111;
        rom_memory[46892] = 3'b111;
        rom_memory[46893] = 3'b110;
        rom_memory[46894] = 3'b110;
        rom_memory[46895] = 3'b110;
        rom_memory[46896] = 3'b110;
        rom_memory[46897] = 3'b110;
        rom_memory[46898] = 3'b110;
        rom_memory[46899] = 3'b110;
        rom_memory[46900] = 3'b110;
        rom_memory[46901] = 3'b110;
        rom_memory[46902] = 3'b110;
        rom_memory[46903] = 3'b111;
        rom_memory[46904] = 3'b111;
        rom_memory[46905] = 3'b111;
        rom_memory[46906] = 3'b111;
        rom_memory[46907] = 3'b111;
        rom_memory[46908] = 3'b111;
        rom_memory[46909] = 3'b111;
        rom_memory[46910] = 3'b111;
        rom_memory[46911] = 3'b111;
        rom_memory[46912] = 3'b111;
        rom_memory[46913] = 3'b111;
        rom_memory[46914] = 3'b111;
        rom_memory[46915] = 3'b111;
        rom_memory[46916] = 3'b111;
        rom_memory[46917] = 3'b110;
        rom_memory[46918] = 3'b110;
        rom_memory[46919] = 3'b110;
        rom_memory[46920] = 3'b110;
        rom_memory[46921] = 3'b110;
        rom_memory[46922] = 3'b110;
        rom_memory[46923] = 3'b110;
        rom_memory[46924] = 3'b110;
        rom_memory[46925] = 3'b110;
        rom_memory[46926] = 3'b110;
        rom_memory[46927] = 3'b110;
        rom_memory[46928] = 3'b110;
        rom_memory[46929] = 3'b110;
        rom_memory[46930] = 3'b110;
        rom_memory[46931] = 3'b110;
        rom_memory[46932] = 3'b110;
        rom_memory[46933] = 3'b110;
        rom_memory[46934] = 3'b110;
        rom_memory[46935] = 3'b110;
        rom_memory[46936] = 3'b110;
        rom_memory[46937] = 3'b110;
        rom_memory[46938] = 3'b110;
        rom_memory[46939] = 3'b110;
        rom_memory[46940] = 3'b110;
        rom_memory[46941] = 3'b110;
        rom_memory[46942] = 3'b110;
        rom_memory[46943] = 3'b110;
        rom_memory[46944] = 3'b110;
        rom_memory[46945] = 3'b110;
        rom_memory[46946] = 3'b110;
        rom_memory[46947] = 3'b110;
        rom_memory[46948] = 3'b110;
        rom_memory[46949] = 3'b110;
        rom_memory[46950] = 3'b110;
        rom_memory[46951] = 3'b110;
        rom_memory[46952] = 3'b110;
        rom_memory[46953] = 3'b110;
        rom_memory[46954] = 3'b110;
        rom_memory[46955] = 3'b110;
        rom_memory[46956] = 3'b110;
        rom_memory[46957] = 3'b110;
        rom_memory[46958] = 3'b110;
        rom_memory[46959] = 3'b110;
        rom_memory[46960] = 3'b110;
        rom_memory[46961] = 3'b110;
        rom_memory[46962] = 3'b110;
        rom_memory[46963] = 3'b110;
        rom_memory[46964] = 3'b110;
        rom_memory[46965] = 3'b110;
        rom_memory[46966] = 3'b110;
        rom_memory[46967] = 3'b110;
        rom_memory[46968] = 3'b110;
        rom_memory[46969] = 3'b110;
        rom_memory[46970] = 3'b110;
        rom_memory[46971] = 3'b110;
        rom_memory[46972] = 3'b110;
        rom_memory[46973] = 3'b110;
        rom_memory[46974] = 3'b110;
        rom_memory[46975] = 3'b110;
        rom_memory[46976] = 3'b110;
        rom_memory[46977] = 3'b110;
        rom_memory[46978] = 3'b110;
        rom_memory[46979] = 3'b110;
        rom_memory[46980] = 3'b110;
        rom_memory[46981] = 3'b110;
        rom_memory[46982] = 3'b110;
        rom_memory[46983] = 3'b110;
        rom_memory[46984] = 3'b110;
        rom_memory[46985] = 3'b110;
        rom_memory[46986] = 3'b110;
        rom_memory[46987] = 3'b110;
        rom_memory[46988] = 3'b110;
        rom_memory[46989] = 3'b110;
        rom_memory[46990] = 3'b110;
        rom_memory[46991] = 3'b110;
        rom_memory[46992] = 3'b110;
        rom_memory[46993] = 3'b110;
        rom_memory[46994] = 3'b110;
        rom_memory[46995] = 3'b110;
        rom_memory[46996] = 3'b110;
        rom_memory[46997] = 3'b110;
        rom_memory[46998] = 3'b110;
        rom_memory[46999] = 3'b110;
        rom_memory[47000] = 3'b110;
        rom_memory[47001] = 3'b110;
        rom_memory[47002] = 3'b110;
        rom_memory[47003] = 3'b110;
        rom_memory[47004] = 3'b110;
        rom_memory[47005] = 3'b110;
        rom_memory[47006] = 3'b110;
        rom_memory[47007] = 3'b110;
        rom_memory[47008] = 3'b110;
        rom_memory[47009] = 3'b110;
        rom_memory[47010] = 3'b110;
        rom_memory[47011] = 3'b110;
        rom_memory[47012] = 3'b110;
        rom_memory[47013] = 3'b110;
        rom_memory[47014] = 3'b110;
        rom_memory[47015] = 3'b110;
        rom_memory[47016] = 3'b110;
        rom_memory[47017] = 3'b110;
        rom_memory[47018] = 3'b100;
        rom_memory[47019] = 3'b000;
        rom_memory[47020] = 3'b000;
        rom_memory[47021] = 3'b000;
        rom_memory[47022] = 3'b000;
        rom_memory[47023] = 3'b000;
        rom_memory[47024] = 3'b100;
        rom_memory[47025] = 3'b110;
        rom_memory[47026] = 3'b110;
        rom_memory[47027] = 3'b110;
        rom_memory[47028] = 3'b110;
        rom_memory[47029] = 3'b110;
        rom_memory[47030] = 3'b110;
        rom_memory[47031] = 3'b110;
        rom_memory[47032] = 3'b110;
        rom_memory[47033] = 3'b110;
        rom_memory[47034] = 3'b110;
        rom_memory[47035] = 3'b110;
        rom_memory[47036] = 3'b110;
        rom_memory[47037] = 3'b110;
        rom_memory[47038] = 3'b110;
        rom_memory[47039] = 3'b110;
        rom_memory[47040] = 3'b111;
        rom_memory[47041] = 3'b111;
        rom_memory[47042] = 3'b111;
        rom_memory[47043] = 3'b111;
        rom_memory[47044] = 3'b111;
        rom_memory[47045] = 3'b111;
        rom_memory[47046] = 3'b111;
        rom_memory[47047] = 3'b111;
        rom_memory[47048] = 3'b111;
        rom_memory[47049] = 3'b111;
        rom_memory[47050] = 3'b111;
        rom_memory[47051] = 3'b111;
        rom_memory[47052] = 3'b111;
        rom_memory[47053] = 3'b111;
        rom_memory[47054] = 3'b111;
        rom_memory[47055] = 3'b111;
        rom_memory[47056] = 3'b110;
        rom_memory[47057] = 3'b110;
        rom_memory[47058] = 3'b110;
        rom_memory[47059] = 3'b110;
        rom_memory[47060] = 3'b110;
        rom_memory[47061] = 3'b110;
        rom_memory[47062] = 3'b110;
        rom_memory[47063] = 3'b110;
        rom_memory[47064] = 3'b110;
        rom_memory[47065] = 3'b110;
        rom_memory[47066] = 3'b110;
        rom_memory[47067] = 3'b110;
        rom_memory[47068] = 3'b110;
        rom_memory[47069] = 3'b110;
        rom_memory[47070] = 3'b110;
        rom_memory[47071] = 3'b110;
        rom_memory[47072] = 3'b110;
        rom_memory[47073] = 3'b111;
        rom_memory[47074] = 3'b111;
        rom_memory[47075] = 3'b111;
        rom_memory[47076] = 3'b111;
        rom_memory[47077] = 3'b111;
        rom_memory[47078] = 3'b110;
        rom_memory[47079] = 3'b110;
        rom_memory[47080] = 3'b110;
        rom_memory[47081] = 3'b110;
        rom_memory[47082] = 3'b111;
        rom_memory[47083] = 3'b111;
        rom_memory[47084] = 3'b111;
        rom_memory[47085] = 3'b110;
        rom_memory[47086] = 3'b110;
        rom_memory[47087] = 3'b111;
        rom_memory[47088] = 3'b111;
        rom_memory[47089] = 3'b111;
        rom_memory[47090] = 3'b110;
        rom_memory[47091] = 3'b110;
        rom_memory[47092] = 3'b110;
        rom_memory[47093] = 3'b110;
        rom_memory[47094] = 3'b110;
        rom_memory[47095] = 3'b110;
        rom_memory[47096] = 3'b111;
        rom_memory[47097] = 3'b110;
        rom_memory[47098] = 3'b110;
        rom_memory[47099] = 3'b110;
        rom_memory[47100] = 3'b110;
        rom_memory[47101] = 3'b100;
        rom_memory[47102] = 3'b100;
        rom_memory[47103] = 3'b110;
        rom_memory[47104] = 3'b110;
        rom_memory[47105] = 3'b110;
        rom_memory[47106] = 3'b000;
        rom_memory[47107] = 3'b100;
        rom_memory[47108] = 3'b111;
        rom_memory[47109] = 3'b111;
        rom_memory[47110] = 3'b111;
        rom_memory[47111] = 3'b111;
        rom_memory[47112] = 3'b110;
        rom_memory[47113] = 3'b111;
        rom_memory[47114] = 3'b111;
        rom_memory[47115] = 3'b000;
        rom_memory[47116] = 3'b000;
        rom_memory[47117] = 3'b111;
        rom_memory[47118] = 3'b111;
        rom_memory[47119] = 3'b000;
        rom_memory[47120] = 3'b100;
        rom_memory[47121] = 3'b110;
        rom_memory[47122] = 3'b110;
        rom_memory[47123] = 3'b110;
        rom_memory[47124] = 3'b110;
        rom_memory[47125] = 3'b110;
        rom_memory[47126] = 3'b110;
        rom_memory[47127] = 3'b111;
        rom_memory[47128] = 3'b111;
        rom_memory[47129] = 3'b110;
        rom_memory[47130] = 3'b110;
        rom_memory[47131] = 3'b111;
        rom_memory[47132] = 3'b111;
        rom_memory[47133] = 3'b110;
        rom_memory[47134] = 3'b110;
        rom_memory[47135] = 3'b110;
        rom_memory[47136] = 3'b110;
        rom_memory[47137] = 3'b110;
        rom_memory[47138] = 3'b110;
        rom_memory[47139] = 3'b110;
        rom_memory[47140] = 3'b110;
        rom_memory[47141] = 3'b110;
        rom_memory[47142] = 3'b110;
        rom_memory[47143] = 3'b110;
        rom_memory[47144] = 3'b111;
        rom_memory[47145] = 3'b111;
        rom_memory[47146] = 3'b111;
        rom_memory[47147] = 3'b111;
        rom_memory[47148] = 3'b111;
        rom_memory[47149] = 3'b111;
        rom_memory[47150] = 3'b111;
        rom_memory[47151] = 3'b111;
        rom_memory[47152] = 3'b111;
        rom_memory[47153] = 3'b111;
        rom_memory[47154] = 3'b111;
        rom_memory[47155] = 3'b111;
        rom_memory[47156] = 3'b111;
        rom_memory[47157] = 3'b110;
        rom_memory[47158] = 3'b110;
        rom_memory[47159] = 3'b110;
        rom_memory[47160] = 3'b110;
        rom_memory[47161] = 3'b110;
        rom_memory[47162] = 3'b110;
        rom_memory[47163] = 3'b110;
        rom_memory[47164] = 3'b110;
        rom_memory[47165] = 3'b110;
        rom_memory[47166] = 3'b110;
        rom_memory[47167] = 3'b110;
        rom_memory[47168] = 3'b110;
        rom_memory[47169] = 3'b110;
        rom_memory[47170] = 3'b110;
        rom_memory[47171] = 3'b110;
        rom_memory[47172] = 3'b110;
        rom_memory[47173] = 3'b110;
        rom_memory[47174] = 3'b110;
        rom_memory[47175] = 3'b110;
        rom_memory[47176] = 3'b110;
        rom_memory[47177] = 3'b110;
        rom_memory[47178] = 3'b110;
        rom_memory[47179] = 3'b110;
        rom_memory[47180] = 3'b110;
        rom_memory[47181] = 3'b110;
        rom_memory[47182] = 3'b110;
        rom_memory[47183] = 3'b110;
        rom_memory[47184] = 3'b110;
        rom_memory[47185] = 3'b110;
        rom_memory[47186] = 3'b110;
        rom_memory[47187] = 3'b110;
        rom_memory[47188] = 3'b110;
        rom_memory[47189] = 3'b110;
        rom_memory[47190] = 3'b110;
        rom_memory[47191] = 3'b110;
        rom_memory[47192] = 3'b110;
        rom_memory[47193] = 3'b110;
        rom_memory[47194] = 3'b110;
        rom_memory[47195] = 3'b110;
        rom_memory[47196] = 3'b110;
        rom_memory[47197] = 3'b110;
        rom_memory[47198] = 3'b110;
        rom_memory[47199] = 3'b110;
        rom_memory[47200] = 3'b110;
        rom_memory[47201] = 3'b110;
        rom_memory[47202] = 3'b110;
        rom_memory[47203] = 3'b110;
        rom_memory[47204] = 3'b110;
        rom_memory[47205] = 3'b110;
        rom_memory[47206] = 3'b110;
        rom_memory[47207] = 3'b110;
        rom_memory[47208] = 3'b110;
        rom_memory[47209] = 3'b110;
        rom_memory[47210] = 3'b110;
        rom_memory[47211] = 3'b110;
        rom_memory[47212] = 3'b110;
        rom_memory[47213] = 3'b110;
        rom_memory[47214] = 3'b110;
        rom_memory[47215] = 3'b110;
        rom_memory[47216] = 3'b110;
        rom_memory[47217] = 3'b110;
        rom_memory[47218] = 3'b110;
        rom_memory[47219] = 3'b110;
        rom_memory[47220] = 3'b110;
        rom_memory[47221] = 3'b110;
        rom_memory[47222] = 3'b110;
        rom_memory[47223] = 3'b110;
        rom_memory[47224] = 3'b110;
        rom_memory[47225] = 3'b110;
        rom_memory[47226] = 3'b110;
        rom_memory[47227] = 3'b110;
        rom_memory[47228] = 3'b110;
        rom_memory[47229] = 3'b110;
        rom_memory[47230] = 3'b110;
        rom_memory[47231] = 3'b110;
        rom_memory[47232] = 3'b110;
        rom_memory[47233] = 3'b110;
        rom_memory[47234] = 3'b110;
        rom_memory[47235] = 3'b110;
        rom_memory[47236] = 3'b110;
        rom_memory[47237] = 3'b110;
        rom_memory[47238] = 3'b110;
        rom_memory[47239] = 3'b110;
        rom_memory[47240] = 3'b110;
        rom_memory[47241] = 3'b110;
        rom_memory[47242] = 3'b110;
        rom_memory[47243] = 3'b110;
        rom_memory[47244] = 3'b110;
        rom_memory[47245] = 3'b110;
        rom_memory[47246] = 3'b110;
        rom_memory[47247] = 3'b110;
        rom_memory[47248] = 3'b110;
        rom_memory[47249] = 3'b110;
        rom_memory[47250] = 3'b110;
        rom_memory[47251] = 3'b110;
        rom_memory[47252] = 3'b110;
        rom_memory[47253] = 3'b110;
        rom_memory[47254] = 3'b110;
        rom_memory[47255] = 3'b110;
        rom_memory[47256] = 3'b110;
        rom_memory[47257] = 3'b110;
        rom_memory[47258] = 3'b110;
        rom_memory[47259] = 3'b110;
        rom_memory[47260] = 3'b000;
        rom_memory[47261] = 3'b000;
        rom_memory[47262] = 3'b000;
        rom_memory[47263] = 3'b000;
        rom_memory[47264] = 3'b000;
        rom_memory[47265] = 3'b000;
        rom_memory[47266] = 3'b110;
        rom_memory[47267] = 3'b110;
        rom_memory[47268] = 3'b110;
        rom_memory[47269] = 3'b110;
        rom_memory[47270] = 3'b110;
        rom_memory[47271] = 3'b110;
        rom_memory[47272] = 3'b110;
        rom_memory[47273] = 3'b110;
        rom_memory[47274] = 3'b110;
        rom_memory[47275] = 3'b110;
        rom_memory[47276] = 3'b110;
        rom_memory[47277] = 3'b110;
        rom_memory[47278] = 3'b110;
        rom_memory[47279] = 3'b110;
        rom_memory[47280] = 3'b110;
        rom_memory[47281] = 3'b111;
        rom_memory[47282] = 3'b111;
        rom_memory[47283] = 3'b111;
        rom_memory[47284] = 3'b111;
        rom_memory[47285] = 3'b111;
        rom_memory[47286] = 3'b111;
        rom_memory[47287] = 3'b111;
        rom_memory[47288] = 3'b111;
        rom_memory[47289] = 3'b111;
        rom_memory[47290] = 3'b111;
        rom_memory[47291] = 3'b111;
        rom_memory[47292] = 3'b111;
        rom_memory[47293] = 3'b111;
        rom_memory[47294] = 3'b111;
        rom_memory[47295] = 3'b111;
        rom_memory[47296] = 3'b110;
        rom_memory[47297] = 3'b110;
        rom_memory[47298] = 3'b110;
        rom_memory[47299] = 3'b110;
        rom_memory[47300] = 3'b110;
        rom_memory[47301] = 3'b110;
        rom_memory[47302] = 3'b110;
        rom_memory[47303] = 3'b110;
        rom_memory[47304] = 3'b110;
        rom_memory[47305] = 3'b110;
        rom_memory[47306] = 3'b110;
        rom_memory[47307] = 3'b110;
        rom_memory[47308] = 3'b110;
        rom_memory[47309] = 3'b110;
        rom_memory[47310] = 3'b110;
        rom_memory[47311] = 3'b110;
        rom_memory[47312] = 3'b110;
        rom_memory[47313] = 3'b110;
        rom_memory[47314] = 3'b110;
        rom_memory[47315] = 3'b111;
        rom_memory[47316] = 3'b111;
        rom_memory[47317] = 3'b110;
        rom_memory[47318] = 3'b110;
        rom_memory[47319] = 3'b110;
        rom_memory[47320] = 3'b110;
        rom_memory[47321] = 3'b110;
        rom_memory[47322] = 3'b111;
        rom_memory[47323] = 3'b111;
        rom_memory[47324] = 3'b111;
        rom_memory[47325] = 3'b110;
        rom_memory[47326] = 3'b110;
        rom_memory[47327] = 3'b110;
        rom_memory[47328] = 3'b111;
        rom_memory[47329] = 3'b111;
        rom_memory[47330] = 3'b110;
        rom_memory[47331] = 3'b110;
        rom_memory[47332] = 3'b110;
        rom_memory[47333] = 3'b110;
        rom_memory[47334] = 3'b110;
        rom_memory[47335] = 3'b110;
        rom_memory[47336] = 3'b111;
        rom_memory[47337] = 3'b110;
        rom_memory[47338] = 3'b110;
        rom_memory[47339] = 3'b110;
        rom_memory[47340] = 3'b110;
        rom_memory[47341] = 3'b110;
        rom_memory[47342] = 3'b100;
        rom_memory[47343] = 3'b100;
        rom_memory[47344] = 3'b100;
        rom_memory[47345] = 3'b110;
        rom_memory[47346] = 3'b000;
        rom_memory[47347] = 3'b000;
        rom_memory[47348] = 3'b111;
        rom_memory[47349] = 3'b111;
        rom_memory[47350] = 3'b100;
        rom_memory[47351] = 3'b111;
        rom_memory[47352] = 3'b111;
        rom_memory[47353] = 3'b000;
        rom_memory[47354] = 3'b000;
        rom_memory[47355] = 3'b111;
        rom_memory[47356] = 3'b111;
        rom_memory[47357] = 3'b111;
        rom_memory[47358] = 3'b111;
        rom_memory[47359] = 3'b111;
        rom_memory[47360] = 3'b111;
        rom_memory[47361] = 3'b111;
        rom_memory[47362] = 3'b110;
        rom_memory[47363] = 3'b100;
        rom_memory[47364] = 3'b100;
        rom_memory[47365] = 3'b110;
        rom_memory[47366] = 3'b110;
        rom_memory[47367] = 3'b110;
        rom_memory[47368] = 3'b110;
        rom_memory[47369] = 3'b110;
        rom_memory[47370] = 3'b111;
        rom_memory[47371] = 3'b110;
        rom_memory[47372] = 3'b110;
        rom_memory[47373] = 3'b110;
        rom_memory[47374] = 3'b110;
        rom_memory[47375] = 3'b110;
        rom_memory[47376] = 3'b110;
        rom_memory[47377] = 3'b110;
        rom_memory[47378] = 3'b110;
        rom_memory[47379] = 3'b110;
        rom_memory[47380] = 3'b110;
        rom_memory[47381] = 3'b110;
        rom_memory[47382] = 3'b110;
        rom_memory[47383] = 3'b110;
        rom_memory[47384] = 3'b110;
        rom_memory[47385] = 3'b111;
        rom_memory[47386] = 3'b111;
        rom_memory[47387] = 3'b111;
        rom_memory[47388] = 3'b111;
        rom_memory[47389] = 3'b111;
        rom_memory[47390] = 3'b111;
        rom_memory[47391] = 3'b111;
        rom_memory[47392] = 3'b111;
        rom_memory[47393] = 3'b111;
        rom_memory[47394] = 3'b111;
        rom_memory[47395] = 3'b111;
        rom_memory[47396] = 3'b111;
        rom_memory[47397] = 3'b111;
        rom_memory[47398] = 3'b110;
        rom_memory[47399] = 3'b110;
        rom_memory[47400] = 3'b110;
        rom_memory[47401] = 3'b110;
        rom_memory[47402] = 3'b110;
        rom_memory[47403] = 3'b110;
        rom_memory[47404] = 3'b110;
        rom_memory[47405] = 3'b110;
        rom_memory[47406] = 3'b110;
        rom_memory[47407] = 3'b110;
        rom_memory[47408] = 3'b110;
        rom_memory[47409] = 3'b110;
        rom_memory[47410] = 3'b110;
        rom_memory[47411] = 3'b110;
        rom_memory[47412] = 3'b110;
        rom_memory[47413] = 3'b110;
        rom_memory[47414] = 3'b110;
        rom_memory[47415] = 3'b110;
        rom_memory[47416] = 3'b110;
        rom_memory[47417] = 3'b110;
        rom_memory[47418] = 3'b110;
        rom_memory[47419] = 3'b110;
        rom_memory[47420] = 3'b110;
        rom_memory[47421] = 3'b110;
        rom_memory[47422] = 3'b110;
        rom_memory[47423] = 3'b110;
        rom_memory[47424] = 3'b110;
        rom_memory[47425] = 3'b110;
        rom_memory[47426] = 3'b110;
        rom_memory[47427] = 3'b110;
        rom_memory[47428] = 3'b110;
        rom_memory[47429] = 3'b110;
        rom_memory[47430] = 3'b110;
        rom_memory[47431] = 3'b110;
        rom_memory[47432] = 3'b110;
        rom_memory[47433] = 3'b110;
        rom_memory[47434] = 3'b110;
        rom_memory[47435] = 3'b110;
        rom_memory[47436] = 3'b110;
        rom_memory[47437] = 3'b110;
        rom_memory[47438] = 3'b110;
        rom_memory[47439] = 3'b110;
        rom_memory[47440] = 3'b110;
        rom_memory[47441] = 3'b110;
        rom_memory[47442] = 3'b110;
        rom_memory[47443] = 3'b110;
        rom_memory[47444] = 3'b110;
        rom_memory[47445] = 3'b110;
        rom_memory[47446] = 3'b110;
        rom_memory[47447] = 3'b110;
        rom_memory[47448] = 3'b110;
        rom_memory[47449] = 3'b110;
        rom_memory[47450] = 3'b110;
        rom_memory[47451] = 3'b110;
        rom_memory[47452] = 3'b110;
        rom_memory[47453] = 3'b110;
        rom_memory[47454] = 3'b110;
        rom_memory[47455] = 3'b110;
        rom_memory[47456] = 3'b110;
        rom_memory[47457] = 3'b110;
        rom_memory[47458] = 3'b110;
        rom_memory[47459] = 3'b110;
        rom_memory[47460] = 3'b110;
        rom_memory[47461] = 3'b110;
        rom_memory[47462] = 3'b110;
        rom_memory[47463] = 3'b110;
        rom_memory[47464] = 3'b110;
        rom_memory[47465] = 3'b110;
        rom_memory[47466] = 3'b110;
        rom_memory[47467] = 3'b110;
        rom_memory[47468] = 3'b110;
        rom_memory[47469] = 3'b110;
        rom_memory[47470] = 3'b110;
        rom_memory[47471] = 3'b110;
        rom_memory[47472] = 3'b110;
        rom_memory[47473] = 3'b110;
        rom_memory[47474] = 3'b110;
        rom_memory[47475] = 3'b110;
        rom_memory[47476] = 3'b110;
        rom_memory[47477] = 3'b110;
        rom_memory[47478] = 3'b110;
        rom_memory[47479] = 3'b110;
        rom_memory[47480] = 3'b110;
        rom_memory[47481] = 3'b110;
        rom_memory[47482] = 3'b110;
        rom_memory[47483] = 3'b110;
        rom_memory[47484] = 3'b110;
        rom_memory[47485] = 3'b110;
        rom_memory[47486] = 3'b110;
        rom_memory[47487] = 3'b110;
        rom_memory[47488] = 3'b110;
        rom_memory[47489] = 3'b110;
        rom_memory[47490] = 3'b110;
        rom_memory[47491] = 3'b110;
        rom_memory[47492] = 3'b110;
        rom_memory[47493] = 3'b110;
        rom_memory[47494] = 3'b110;
        rom_memory[47495] = 3'b110;
        rom_memory[47496] = 3'b110;
        rom_memory[47497] = 3'b110;
        rom_memory[47498] = 3'b110;
        rom_memory[47499] = 3'b110;
        rom_memory[47500] = 3'b110;
        rom_memory[47501] = 3'b110;
        rom_memory[47502] = 3'b100;
        rom_memory[47503] = 3'b000;
        rom_memory[47504] = 3'b000;
        rom_memory[47505] = 3'b000;
        rom_memory[47506] = 3'b000;
        rom_memory[47507] = 3'b100;
        rom_memory[47508] = 3'b110;
        rom_memory[47509] = 3'b110;
        rom_memory[47510] = 3'b110;
        rom_memory[47511] = 3'b110;
        rom_memory[47512] = 3'b110;
        rom_memory[47513] = 3'b110;
        rom_memory[47514] = 3'b110;
        rom_memory[47515] = 3'b110;
        rom_memory[47516] = 3'b110;
        rom_memory[47517] = 3'b110;
        rom_memory[47518] = 3'b110;
        rom_memory[47519] = 3'b110;
        rom_memory[47520] = 3'b110;
        rom_memory[47521] = 3'b111;
        rom_memory[47522] = 3'b111;
        rom_memory[47523] = 3'b111;
        rom_memory[47524] = 3'b111;
        rom_memory[47525] = 3'b111;
        rom_memory[47526] = 3'b111;
        rom_memory[47527] = 3'b111;
        rom_memory[47528] = 3'b111;
        rom_memory[47529] = 3'b111;
        rom_memory[47530] = 3'b111;
        rom_memory[47531] = 3'b111;
        rom_memory[47532] = 3'b111;
        rom_memory[47533] = 3'b111;
        rom_memory[47534] = 3'b111;
        rom_memory[47535] = 3'b110;
        rom_memory[47536] = 3'b110;
        rom_memory[47537] = 3'b110;
        rom_memory[47538] = 3'b110;
        rom_memory[47539] = 3'b110;
        rom_memory[47540] = 3'b110;
        rom_memory[47541] = 3'b110;
        rom_memory[47542] = 3'b110;
        rom_memory[47543] = 3'b110;
        rom_memory[47544] = 3'b110;
        rom_memory[47545] = 3'b110;
        rom_memory[47546] = 3'b110;
        rom_memory[47547] = 3'b110;
        rom_memory[47548] = 3'b110;
        rom_memory[47549] = 3'b110;
        rom_memory[47550] = 3'b110;
        rom_memory[47551] = 3'b110;
        rom_memory[47552] = 3'b110;
        rom_memory[47553] = 3'b110;
        rom_memory[47554] = 3'b110;
        rom_memory[47555] = 3'b111;
        rom_memory[47556] = 3'b110;
        rom_memory[47557] = 3'b110;
        rom_memory[47558] = 3'b110;
        rom_memory[47559] = 3'b110;
        rom_memory[47560] = 3'b110;
        rom_memory[47561] = 3'b110;
        rom_memory[47562] = 3'b111;
        rom_memory[47563] = 3'b111;
        rom_memory[47564] = 3'b111;
        rom_memory[47565] = 3'b110;
        rom_memory[47566] = 3'b110;
        rom_memory[47567] = 3'b110;
        rom_memory[47568] = 3'b111;
        rom_memory[47569] = 3'b111;
        rom_memory[47570] = 3'b110;
        rom_memory[47571] = 3'b110;
        rom_memory[47572] = 3'b110;
        rom_memory[47573] = 3'b110;
        rom_memory[47574] = 3'b110;
        rom_memory[47575] = 3'b111;
        rom_memory[47576] = 3'b111;
        rom_memory[47577] = 3'b110;
        rom_memory[47578] = 3'b110;
        rom_memory[47579] = 3'b110;
        rom_memory[47580] = 3'b110;
        rom_memory[47581] = 3'b110;
        rom_memory[47582] = 3'b110;
        rom_memory[47583] = 3'b110;
        rom_memory[47584] = 3'b111;
        rom_memory[47585] = 3'b111;
        rom_memory[47586] = 3'b111;
        rom_memory[47587] = 3'b000;
        rom_memory[47588] = 3'b111;
        rom_memory[47589] = 3'b111;
        rom_memory[47590] = 3'b000;
        rom_memory[47591] = 3'b100;
        rom_memory[47592] = 3'b100;
        rom_memory[47593] = 3'b000;
        rom_memory[47594] = 3'b111;
        rom_memory[47595] = 3'b111;
        rom_memory[47596] = 3'b111;
        rom_memory[47597] = 3'b111;
        rom_memory[47598] = 3'b111;
        rom_memory[47599] = 3'b111;
        rom_memory[47600] = 3'b111;
        rom_memory[47601] = 3'b111;
        rom_memory[47602] = 3'b111;
        rom_memory[47603] = 3'b100;
        rom_memory[47604] = 3'b110;
        rom_memory[47605] = 3'b110;
        rom_memory[47606] = 3'b110;
        rom_memory[47607] = 3'b110;
        rom_memory[47608] = 3'b110;
        rom_memory[47609] = 3'b111;
        rom_memory[47610] = 3'b110;
        rom_memory[47611] = 3'b110;
        rom_memory[47612] = 3'b110;
        rom_memory[47613] = 3'b110;
        rom_memory[47614] = 3'b110;
        rom_memory[47615] = 3'b110;
        rom_memory[47616] = 3'b110;
        rom_memory[47617] = 3'b110;
        rom_memory[47618] = 3'b110;
        rom_memory[47619] = 3'b110;
        rom_memory[47620] = 3'b110;
        rom_memory[47621] = 3'b100;
        rom_memory[47622] = 3'b100;
        rom_memory[47623] = 3'b100;
        rom_memory[47624] = 3'b110;
        rom_memory[47625] = 3'b110;
        rom_memory[47626] = 3'b110;
        rom_memory[47627] = 3'b111;
        rom_memory[47628] = 3'b111;
        rom_memory[47629] = 3'b111;
        rom_memory[47630] = 3'b111;
        rom_memory[47631] = 3'b111;
        rom_memory[47632] = 3'b111;
        rom_memory[47633] = 3'b111;
        rom_memory[47634] = 3'b111;
        rom_memory[47635] = 3'b111;
        rom_memory[47636] = 3'b111;
        rom_memory[47637] = 3'b111;
        rom_memory[47638] = 3'b110;
        rom_memory[47639] = 3'b110;
        rom_memory[47640] = 3'b110;
        rom_memory[47641] = 3'b110;
        rom_memory[47642] = 3'b110;
        rom_memory[47643] = 3'b110;
        rom_memory[47644] = 3'b110;
        rom_memory[47645] = 3'b110;
        rom_memory[47646] = 3'b110;
        rom_memory[47647] = 3'b110;
        rom_memory[47648] = 3'b110;
        rom_memory[47649] = 3'b110;
        rom_memory[47650] = 3'b110;
        rom_memory[47651] = 3'b110;
        rom_memory[47652] = 3'b110;
        rom_memory[47653] = 3'b110;
        rom_memory[47654] = 3'b110;
        rom_memory[47655] = 3'b110;
        rom_memory[47656] = 3'b110;
        rom_memory[47657] = 3'b110;
        rom_memory[47658] = 3'b110;
        rom_memory[47659] = 3'b110;
        rom_memory[47660] = 3'b110;
        rom_memory[47661] = 3'b110;
        rom_memory[47662] = 3'b110;
        rom_memory[47663] = 3'b110;
        rom_memory[47664] = 3'b110;
        rom_memory[47665] = 3'b110;
        rom_memory[47666] = 3'b110;
        rom_memory[47667] = 3'b110;
        rom_memory[47668] = 3'b110;
        rom_memory[47669] = 3'b110;
        rom_memory[47670] = 3'b110;
        rom_memory[47671] = 3'b110;
        rom_memory[47672] = 3'b110;
        rom_memory[47673] = 3'b110;
        rom_memory[47674] = 3'b110;
        rom_memory[47675] = 3'b110;
        rom_memory[47676] = 3'b110;
        rom_memory[47677] = 3'b110;
        rom_memory[47678] = 3'b110;
        rom_memory[47679] = 3'b110;
        rom_memory[47680] = 3'b110;
        rom_memory[47681] = 3'b110;
        rom_memory[47682] = 3'b110;
        rom_memory[47683] = 3'b110;
        rom_memory[47684] = 3'b110;
        rom_memory[47685] = 3'b110;
        rom_memory[47686] = 3'b110;
        rom_memory[47687] = 3'b110;
        rom_memory[47688] = 3'b110;
        rom_memory[47689] = 3'b110;
        rom_memory[47690] = 3'b110;
        rom_memory[47691] = 3'b110;
        rom_memory[47692] = 3'b110;
        rom_memory[47693] = 3'b110;
        rom_memory[47694] = 3'b110;
        rom_memory[47695] = 3'b110;
        rom_memory[47696] = 3'b110;
        rom_memory[47697] = 3'b110;
        rom_memory[47698] = 3'b110;
        rom_memory[47699] = 3'b110;
        rom_memory[47700] = 3'b110;
        rom_memory[47701] = 3'b110;
        rom_memory[47702] = 3'b110;
        rom_memory[47703] = 3'b110;
        rom_memory[47704] = 3'b110;
        rom_memory[47705] = 3'b110;
        rom_memory[47706] = 3'b110;
        rom_memory[47707] = 3'b110;
        rom_memory[47708] = 3'b110;
        rom_memory[47709] = 3'b110;
        rom_memory[47710] = 3'b110;
        rom_memory[47711] = 3'b110;
        rom_memory[47712] = 3'b110;
        rom_memory[47713] = 3'b110;
        rom_memory[47714] = 3'b110;
        rom_memory[47715] = 3'b110;
        rom_memory[47716] = 3'b110;
        rom_memory[47717] = 3'b110;
        rom_memory[47718] = 3'b110;
        rom_memory[47719] = 3'b110;
        rom_memory[47720] = 3'b110;
        rom_memory[47721] = 3'b110;
        rom_memory[47722] = 3'b110;
        rom_memory[47723] = 3'b110;
        rom_memory[47724] = 3'b110;
        rom_memory[47725] = 3'b110;
        rom_memory[47726] = 3'b110;
        rom_memory[47727] = 3'b110;
        rom_memory[47728] = 3'b110;
        rom_memory[47729] = 3'b110;
        rom_memory[47730] = 3'b110;
        rom_memory[47731] = 3'b110;
        rom_memory[47732] = 3'b110;
        rom_memory[47733] = 3'b110;
        rom_memory[47734] = 3'b110;
        rom_memory[47735] = 3'b110;
        rom_memory[47736] = 3'b110;
        rom_memory[47737] = 3'b110;
        rom_memory[47738] = 3'b110;
        rom_memory[47739] = 3'b110;
        rom_memory[47740] = 3'b110;
        rom_memory[47741] = 3'b110;
        rom_memory[47742] = 3'b110;
        rom_memory[47743] = 3'b110;
        rom_memory[47744] = 3'b110;
        rom_memory[47745] = 3'b110;
        rom_memory[47746] = 3'b000;
        rom_memory[47747] = 3'b100;
        rom_memory[47748] = 3'b110;
        rom_memory[47749] = 3'b110;
        rom_memory[47750] = 3'b110;
        rom_memory[47751] = 3'b110;
        rom_memory[47752] = 3'b110;
        rom_memory[47753] = 3'b110;
        rom_memory[47754] = 3'b110;
        rom_memory[47755] = 3'b110;
        rom_memory[47756] = 3'b110;
        rom_memory[47757] = 3'b110;
        rom_memory[47758] = 3'b110;
        rom_memory[47759] = 3'b110;
        rom_memory[47760] = 3'b110;
        rom_memory[47761] = 3'b111;
        rom_memory[47762] = 3'b111;
        rom_memory[47763] = 3'b111;
        rom_memory[47764] = 3'b111;
        rom_memory[47765] = 3'b111;
        rom_memory[47766] = 3'b111;
        rom_memory[47767] = 3'b111;
        rom_memory[47768] = 3'b111;
        rom_memory[47769] = 3'b111;
        rom_memory[47770] = 3'b111;
        rom_memory[47771] = 3'b111;
        rom_memory[47772] = 3'b111;
        rom_memory[47773] = 3'b111;
        rom_memory[47774] = 3'b111;
        rom_memory[47775] = 3'b110;
        rom_memory[47776] = 3'b110;
        rom_memory[47777] = 3'b110;
        rom_memory[47778] = 3'b110;
        rom_memory[47779] = 3'b110;
        rom_memory[47780] = 3'b110;
        rom_memory[47781] = 3'b110;
        rom_memory[47782] = 3'b110;
        rom_memory[47783] = 3'b110;
        rom_memory[47784] = 3'b110;
        rom_memory[47785] = 3'b110;
        rom_memory[47786] = 3'b110;
        rom_memory[47787] = 3'b110;
        rom_memory[47788] = 3'b110;
        rom_memory[47789] = 3'b110;
        rom_memory[47790] = 3'b110;
        rom_memory[47791] = 3'b110;
        rom_memory[47792] = 3'b110;
        rom_memory[47793] = 3'b110;
        rom_memory[47794] = 3'b110;
        rom_memory[47795] = 3'b110;
        rom_memory[47796] = 3'b110;
        rom_memory[47797] = 3'b110;
        rom_memory[47798] = 3'b110;
        rom_memory[47799] = 3'b110;
        rom_memory[47800] = 3'b110;
        rom_memory[47801] = 3'b110;
        rom_memory[47802] = 3'b110;
        rom_memory[47803] = 3'b111;
        rom_memory[47804] = 3'b111;
        rom_memory[47805] = 3'b110;
        rom_memory[47806] = 3'b110;
        rom_memory[47807] = 3'b110;
        rom_memory[47808] = 3'b110;
        rom_memory[47809] = 3'b110;
        rom_memory[47810] = 3'b110;
        rom_memory[47811] = 3'b110;
        rom_memory[47812] = 3'b110;
        rom_memory[47813] = 3'b110;
        rom_memory[47814] = 3'b110;
        rom_memory[47815] = 3'b111;
        rom_memory[47816] = 3'b111;
        rom_memory[47817] = 3'b110;
        rom_memory[47818] = 3'b110;
        rom_memory[47819] = 3'b110;
        rom_memory[47820] = 3'b110;
        rom_memory[47821] = 3'b110;
        rom_memory[47822] = 3'b110;
        rom_memory[47823] = 3'b111;
        rom_memory[47824] = 3'b111;
        rom_memory[47825] = 3'b111;
        rom_memory[47826] = 3'b110;
        rom_memory[47827] = 3'b000;
        rom_memory[47828] = 3'b000;
        rom_memory[47829] = 3'b111;
        rom_memory[47830] = 3'b000;
        rom_memory[47831] = 3'b111;
        rom_memory[47832] = 3'b100;
        rom_memory[47833] = 3'b000;
        rom_memory[47834] = 3'b111;
        rom_memory[47835] = 3'b111;
        rom_memory[47836] = 3'b111;
        rom_memory[47837] = 3'b111;
        rom_memory[47838] = 3'b111;
        rom_memory[47839] = 3'b111;
        rom_memory[47840] = 3'b111;
        rom_memory[47841] = 3'b111;
        rom_memory[47842] = 3'b111;
        rom_memory[47843] = 3'b110;
        rom_memory[47844] = 3'b110;
        rom_memory[47845] = 3'b110;
        rom_memory[47846] = 3'b110;
        rom_memory[47847] = 3'b110;
        rom_memory[47848] = 3'b110;
        rom_memory[47849] = 3'b111;
        rom_memory[47850] = 3'b110;
        rom_memory[47851] = 3'b110;
        rom_memory[47852] = 3'b110;
        rom_memory[47853] = 3'b110;
        rom_memory[47854] = 3'b110;
        rom_memory[47855] = 3'b110;
        rom_memory[47856] = 3'b110;
        rom_memory[47857] = 3'b110;
        rom_memory[47858] = 3'b110;
        rom_memory[47859] = 3'b110;
        rom_memory[47860] = 3'b110;
        rom_memory[47861] = 3'b110;
        rom_memory[47862] = 3'b100;
        rom_memory[47863] = 3'b100;
        rom_memory[47864] = 3'b100;
        rom_memory[47865] = 3'b100;
        rom_memory[47866] = 3'b100;
        rom_memory[47867] = 3'b100;
        rom_memory[47868] = 3'b111;
        rom_memory[47869] = 3'b111;
        rom_memory[47870] = 3'b111;
        rom_memory[47871] = 3'b111;
        rom_memory[47872] = 3'b111;
        rom_memory[47873] = 3'b111;
        rom_memory[47874] = 3'b110;
        rom_memory[47875] = 3'b110;
        rom_memory[47876] = 3'b111;
        rom_memory[47877] = 3'b111;
        rom_memory[47878] = 3'b111;
        rom_memory[47879] = 3'b110;
        rom_memory[47880] = 3'b110;
        rom_memory[47881] = 3'b110;
        rom_memory[47882] = 3'b110;
        rom_memory[47883] = 3'b110;
        rom_memory[47884] = 3'b110;
        rom_memory[47885] = 3'b110;
        rom_memory[47886] = 3'b110;
        rom_memory[47887] = 3'b110;
        rom_memory[47888] = 3'b110;
        rom_memory[47889] = 3'b110;
        rom_memory[47890] = 3'b110;
        rom_memory[47891] = 3'b110;
        rom_memory[47892] = 3'b110;
        rom_memory[47893] = 3'b110;
        rom_memory[47894] = 3'b110;
        rom_memory[47895] = 3'b110;
        rom_memory[47896] = 3'b110;
        rom_memory[47897] = 3'b110;
        rom_memory[47898] = 3'b110;
        rom_memory[47899] = 3'b110;
        rom_memory[47900] = 3'b110;
        rom_memory[47901] = 3'b110;
        rom_memory[47902] = 3'b110;
        rom_memory[47903] = 3'b110;
        rom_memory[47904] = 3'b110;
        rom_memory[47905] = 3'b110;
        rom_memory[47906] = 3'b110;
        rom_memory[47907] = 3'b110;
        rom_memory[47908] = 3'b110;
        rom_memory[47909] = 3'b110;
        rom_memory[47910] = 3'b110;
        rom_memory[47911] = 3'b110;
        rom_memory[47912] = 3'b110;
        rom_memory[47913] = 3'b110;
        rom_memory[47914] = 3'b110;
        rom_memory[47915] = 3'b110;
        rom_memory[47916] = 3'b110;
        rom_memory[47917] = 3'b110;
        rom_memory[47918] = 3'b110;
        rom_memory[47919] = 3'b110;
        rom_memory[47920] = 3'b110;
        rom_memory[47921] = 3'b110;
        rom_memory[47922] = 3'b110;
        rom_memory[47923] = 3'b110;
        rom_memory[47924] = 3'b110;
        rom_memory[47925] = 3'b110;
        rom_memory[47926] = 3'b110;
        rom_memory[47927] = 3'b110;
        rom_memory[47928] = 3'b110;
        rom_memory[47929] = 3'b110;
        rom_memory[47930] = 3'b110;
        rom_memory[47931] = 3'b110;
        rom_memory[47932] = 3'b110;
        rom_memory[47933] = 3'b110;
        rom_memory[47934] = 3'b110;
        rom_memory[47935] = 3'b110;
        rom_memory[47936] = 3'b110;
        rom_memory[47937] = 3'b110;
        rom_memory[47938] = 3'b110;
        rom_memory[47939] = 3'b110;
        rom_memory[47940] = 3'b110;
        rom_memory[47941] = 3'b110;
        rom_memory[47942] = 3'b110;
        rom_memory[47943] = 3'b110;
        rom_memory[47944] = 3'b110;
        rom_memory[47945] = 3'b110;
        rom_memory[47946] = 3'b110;
        rom_memory[47947] = 3'b110;
        rom_memory[47948] = 3'b110;
        rom_memory[47949] = 3'b110;
        rom_memory[47950] = 3'b110;
        rom_memory[47951] = 3'b110;
        rom_memory[47952] = 3'b110;
        rom_memory[47953] = 3'b110;
        rom_memory[47954] = 3'b110;
        rom_memory[47955] = 3'b110;
        rom_memory[47956] = 3'b110;
        rom_memory[47957] = 3'b110;
        rom_memory[47958] = 3'b110;
        rom_memory[47959] = 3'b110;
        rom_memory[47960] = 3'b110;
        rom_memory[47961] = 3'b110;
        rom_memory[47962] = 3'b110;
        rom_memory[47963] = 3'b110;
        rom_memory[47964] = 3'b110;
        rom_memory[47965] = 3'b110;
        rom_memory[47966] = 3'b110;
        rom_memory[47967] = 3'b110;
        rom_memory[47968] = 3'b110;
        rom_memory[47969] = 3'b110;
        rom_memory[47970] = 3'b110;
        rom_memory[47971] = 3'b110;
        rom_memory[47972] = 3'b110;
        rom_memory[47973] = 3'b110;
        rom_memory[47974] = 3'b110;
        rom_memory[47975] = 3'b110;
        rom_memory[47976] = 3'b110;
        rom_memory[47977] = 3'b110;
        rom_memory[47978] = 3'b110;
        rom_memory[47979] = 3'b110;
        rom_memory[47980] = 3'b110;
        rom_memory[47981] = 3'b110;
        rom_memory[47982] = 3'b110;
        rom_memory[47983] = 3'b110;
        rom_memory[47984] = 3'b110;
        rom_memory[47985] = 3'b110;
        rom_memory[47986] = 3'b110;
        rom_memory[47987] = 3'b110;
        rom_memory[47988] = 3'b110;
        rom_memory[47989] = 3'b110;
        rom_memory[47990] = 3'b110;
        rom_memory[47991] = 3'b110;
        rom_memory[47992] = 3'b110;
        rom_memory[47993] = 3'b110;
        rom_memory[47994] = 3'b110;
        rom_memory[47995] = 3'b110;
        rom_memory[47996] = 3'b110;
        rom_memory[47997] = 3'b110;
        rom_memory[47998] = 3'b110;
        rom_memory[47999] = 3'b110;
        rom_memory[48000] = 3'b110;
        rom_memory[48001] = 3'b111;
        rom_memory[48002] = 3'b111;
        rom_memory[48003] = 3'b111;
        rom_memory[48004] = 3'b110;
        rom_memory[48005] = 3'b111;
        rom_memory[48006] = 3'b111;
        rom_memory[48007] = 3'b111;
        rom_memory[48008] = 3'b111;
        rom_memory[48009] = 3'b111;
        rom_memory[48010] = 3'b111;
        rom_memory[48011] = 3'b111;
        rom_memory[48012] = 3'b111;
        rom_memory[48013] = 3'b111;
        rom_memory[48014] = 3'b111;
        rom_memory[48015] = 3'b110;
        rom_memory[48016] = 3'b110;
        rom_memory[48017] = 3'b110;
        rom_memory[48018] = 3'b110;
        rom_memory[48019] = 3'b110;
        rom_memory[48020] = 3'b110;
        rom_memory[48021] = 3'b110;
        rom_memory[48022] = 3'b110;
        rom_memory[48023] = 3'b110;
        rom_memory[48024] = 3'b110;
        rom_memory[48025] = 3'b110;
        rom_memory[48026] = 3'b110;
        rom_memory[48027] = 3'b110;
        rom_memory[48028] = 3'b110;
        rom_memory[48029] = 3'b110;
        rom_memory[48030] = 3'b110;
        rom_memory[48031] = 3'b110;
        rom_memory[48032] = 3'b110;
        rom_memory[48033] = 3'b110;
        rom_memory[48034] = 3'b110;
        rom_memory[48035] = 3'b110;
        rom_memory[48036] = 3'b110;
        rom_memory[48037] = 3'b110;
        rom_memory[48038] = 3'b110;
        rom_memory[48039] = 3'b110;
        rom_memory[48040] = 3'b110;
        rom_memory[48041] = 3'b110;
        rom_memory[48042] = 3'b110;
        rom_memory[48043] = 3'b111;
        rom_memory[48044] = 3'b111;
        rom_memory[48045] = 3'b111;
        rom_memory[48046] = 3'b110;
        rom_memory[48047] = 3'b110;
        rom_memory[48048] = 3'b110;
        rom_memory[48049] = 3'b110;
        rom_memory[48050] = 3'b111;
        rom_memory[48051] = 3'b110;
        rom_memory[48052] = 3'b110;
        rom_memory[48053] = 3'b110;
        rom_memory[48054] = 3'b110;
        rom_memory[48055] = 3'b111;
        rom_memory[48056] = 3'b111;
        rom_memory[48057] = 3'b111;
        rom_memory[48058] = 3'b110;
        rom_memory[48059] = 3'b110;
        rom_memory[48060] = 3'b110;
        rom_memory[48061] = 3'b111;
        rom_memory[48062] = 3'b111;
        rom_memory[48063] = 3'b111;
        rom_memory[48064] = 3'b111;
        rom_memory[48065] = 3'b111;
        rom_memory[48066] = 3'b111;
        rom_memory[48067] = 3'b100;
        rom_memory[48068] = 3'b000;
        rom_memory[48069] = 3'b000;
        rom_memory[48070] = 3'b111;
        rom_memory[48071] = 3'b111;
        rom_memory[48072] = 3'b111;
        rom_memory[48073] = 3'b100;
        rom_memory[48074] = 3'b111;
        rom_memory[48075] = 3'b111;
        rom_memory[48076] = 3'b111;
        rom_memory[48077] = 3'b111;
        rom_memory[48078] = 3'b111;
        rom_memory[48079] = 3'b111;
        rom_memory[48080] = 3'b111;
        rom_memory[48081] = 3'b111;
        rom_memory[48082] = 3'b110;
        rom_memory[48083] = 3'b100;
        rom_memory[48084] = 3'b100;
        rom_memory[48085] = 3'b100;
        rom_memory[48086] = 3'b110;
        rom_memory[48087] = 3'b110;
        rom_memory[48088] = 3'b111;
        rom_memory[48089] = 3'b111;
        rom_memory[48090] = 3'b110;
        rom_memory[48091] = 3'b110;
        rom_memory[48092] = 3'b110;
        rom_memory[48093] = 3'b110;
        rom_memory[48094] = 3'b110;
        rom_memory[48095] = 3'b110;
        rom_memory[48096] = 3'b110;
        rom_memory[48097] = 3'b110;
        rom_memory[48098] = 3'b110;
        rom_memory[48099] = 3'b110;
        rom_memory[48100] = 3'b110;
        rom_memory[48101] = 3'b110;
        rom_memory[48102] = 3'b110;
        rom_memory[48103] = 3'b100;
        rom_memory[48104] = 3'b000;
        rom_memory[48105] = 3'b000;
        rom_memory[48106] = 3'b000;
        rom_memory[48107] = 3'b100;
        rom_memory[48108] = 3'b100;
        rom_memory[48109] = 3'b111;
        rom_memory[48110] = 3'b111;
        rom_memory[48111] = 3'b111;
        rom_memory[48112] = 3'b111;
        rom_memory[48113] = 3'b111;
        rom_memory[48114] = 3'b100;
        rom_memory[48115] = 3'b111;
        rom_memory[48116] = 3'b111;
        rom_memory[48117] = 3'b111;
        rom_memory[48118] = 3'b111;
        rom_memory[48119] = 3'b111;
        rom_memory[48120] = 3'b110;
        rom_memory[48121] = 3'b110;
        rom_memory[48122] = 3'b110;
        rom_memory[48123] = 3'b110;
        rom_memory[48124] = 3'b110;
        rom_memory[48125] = 3'b110;
        rom_memory[48126] = 3'b110;
        rom_memory[48127] = 3'b110;
        rom_memory[48128] = 3'b110;
        rom_memory[48129] = 3'b110;
        rom_memory[48130] = 3'b110;
        rom_memory[48131] = 3'b110;
        rom_memory[48132] = 3'b110;
        rom_memory[48133] = 3'b110;
        rom_memory[48134] = 3'b110;
        rom_memory[48135] = 3'b110;
        rom_memory[48136] = 3'b110;
        rom_memory[48137] = 3'b110;
        rom_memory[48138] = 3'b110;
        rom_memory[48139] = 3'b110;
        rom_memory[48140] = 3'b110;
        rom_memory[48141] = 3'b110;
        rom_memory[48142] = 3'b110;
        rom_memory[48143] = 3'b110;
        rom_memory[48144] = 3'b110;
        rom_memory[48145] = 3'b110;
        rom_memory[48146] = 3'b110;
        rom_memory[48147] = 3'b110;
        rom_memory[48148] = 3'b110;
        rom_memory[48149] = 3'b110;
        rom_memory[48150] = 3'b110;
        rom_memory[48151] = 3'b110;
        rom_memory[48152] = 3'b110;
        rom_memory[48153] = 3'b110;
        rom_memory[48154] = 3'b110;
        rom_memory[48155] = 3'b110;
        rom_memory[48156] = 3'b110;
        rom_memory[48157] = 3'b110;
        rom_memory[48158] = 3'b110;
        rom_memory[48159] = 3'b110;
        rom_memory[48160] = 3'b110;
        rom_memory[48161] = 3'b110;
        rom_memory[48162] = 3'b110;
        rom_memory[48163] = 3'b110;
        rom_memory[48164] = 3'b110;
        rom_memory[48165] = 3'b110;
        rom_memory[48166] = 3'b110;
        rom_memory[48167] = 3'b110;
        rom_memory[48168] = 3'b110;
        rom_memory[48169] = 3'b110;
        rom_memory[48170] = 3'b110;
        rom_memory[48171] = 3'b110;
        rom_memory[48172] = 3'b110;
        rom_memory[48173] = 3'b110;
        rom_memory[48174] = 3'b110;
        rom_memory[48175] = 3'b110;
        rom_memory[48176] = 3'b110;
        rom_memory[48177] = 3'b110;
        rom_memory[48178] = 3'b110;
        rom_memory[48179] = 3'b110;
        rom_memory[48180] = 3'b110;
        rom_memory[48181] = 3'b110;
        rom_memory[48182] = 3'b110;
        rom_memory[48183] = 3'b110;
        rom_memory[48184] = 3'b110;
        rom_memory[48185] = 3'b110;
        rom_memory[48186] = 3'b110;
        rom_memory[48187] = 3'b110;
        rom_memory[48188] = 3'b110;
        rom_memory[48189] = 3'b110;
        rom_memory[48190] = 3'b110;
        rom_memory[48191] = 3'b110;
        rom_memory[48192] = 3'b110;
        rom_memory[48193] = 3'b110;
        rom_memory[48194] = 3'b110;
        rom_memory[48195] = 3'b110;
        rom_memory[48196] = 3'b110;
        rom_memory[48197] = 3'b110;
        rom_memory[48198] = 3'b110;
        rom_memory[48199] = 3'b110;
        rom_memory[48200] = 3'b110;
        rom_memory[48201] = 3'b110;
        rom_memory[48202] = 3'b110;
        rom_memory[48203] = 3'b110;
        rom_memory[48204] = 3'b110;
        rom_memory[48205] = 3'b110;
        rom_memory[48206] = 3'b110;
        rom_memory[48207] = 3'b110;
        rom_memory[48208] = 3'b110;
        rom_memory[48209] = 3'b110;
        rom_memory[48210] = 3'b110;
        rom_memory[48211] = 3'b110;
        rom_memory[48212] = 3'b110;
        rom_memory[48213] = 3'b110;
        rom_memory[48214] = 3'b110;
        rom_memory[48215] = 3'b110;
        rom_memory[48216] = 3'b110;
        rom_memory[48217] = 3'b110;
        rom_memory[48218] = 3'b110;
        rom_memory[48219] = 3'b110;
        rom_memory[48220] = 3'b110;
        rom_memory[48221] = 3'b110;
        rom_memory[48222] = 3'b110;
        rom_memory[48223] = 3'b110;
        rom_memory[48224] = 3'b110;
        rom_memory[48225] = 3'b110;
        rom_memory[48226] = 3'b110;
        rom_memory[48227] = 3'b110;
        rom_memory[48228] = 3'b110;
        rom_memory[48229] = 3'b110;
        rom_memory[48230] = 3'b110;
        rom_memory[48231] = 3'b110;
        rom_memory[48232] = 3'b110;
        rom_memory[48233] = 3'b110;
        rom_memory[48234] = 3'b110;
        rom_memory[48235] = 3'b110;
        rom_memory[48236] = 3'b110;
        rom_memory[48237] = 3'b110;
        rom_memory[48238] = 3'b110;
        rom_memory[48239] = 3'b110;
        rom_memory[48240] = 3'b110;
        rom_memory[48241] = 3'b110;
        rom_memory[48242] = 3'b111;
        rom_memory[48243] = 3'b111;
        rom_memory[48244] = 3'b110;
        rom_memory[48245] = 3'b111;
        rom_memory[48246] = 3'b111;
        rom_memory[48247] = 3'b111;
        rom_memory[48248] = 3'b111;
        rom_memory[48249] = 3'b111;
        rom_memory[48250] = 3'b111;
        rom_memory[48251] = 3'b111;
        rom_memory[48252] = 3'b111;
        rom_memory[48253] = 3'b111;
        rom_memory[48254] = 3'b110;
        rom_memory[48255] = 3'b110;
        rom_memory[48256] = 3'b110;
        rom_memory[48257] = 3'b110;
        rom_memory[48258] = 3'b110;
        rom_memory[48259] = 3'b110;
        rom_memory[48260] = 3'b110;
        rom_memory[48261] = 3'b110;
        rom_memory[48262] = 3'b110;
        rom_memory[48263] = 3'b110;
        rom_memory[48264] = 3'b110;
        rom_memory[48265] = 3'b110;
        rom_memory[48266] = 3'b110;
        rom_memory[48267] = 3'b110;
        rom_memory[48268] = 3'b110;
        rom_memory[48269] = 3'b110;
        rom_memory[48270] = 3'b110;
        rom_memory[48271] = 3'b110;
        rom_memory[48272] = 3'b110;
        rom_memory[48273] = 3'b110;
        rom_memory[48274] = 3'b110;
        rom_memory[48275] = 3'b110;
        rom_memory[48276] = 3'b110;
        rom_memory[48277] = 3'b110;
        rom_memory[48278] = 3'b110;
        rom_memory[48279] = 3'b110;
        rom_memory[48280] = 3'b110;
        rom_memory[48281] = 3'b110;
        rom_memory[48282] = 3'b110;
        rom_memory[48283] = 3'b110;
        rom_memory[48284] = 3'b111;
        rom_memory[48285] = 3'b111;
        rom_memory[48286] = 3'b110;
        rom_memory[48287] = 3'b110;
        rom_memory[48288] = 3'b110;
        rom_memory[48289] = 3'b110;
        rom_memory[48290] = 3'b110;
        rom_memory[48291] = 3'b110;
        rom_memory[48292] = 3'b110;
        rom_memory[48293] = 3'b111;
        rom_memory[48294] = 3'b111;
        rom_memory[48295] = 3'b111;
        rom_memory[48296] = 3'b111;
        rom_memory[48297] = 3'b111;
        rom_memory[48298] = 3'b111;
        rom_memory[48299] = 3'b111;
        rom_memory[48300] = 3'b111;
        rom_memory[48301] = 3'b111;
        rom_memory[48302] = 3'b111;
        rom_memory[48303] = 3'b110;
        rom_memory[48304] = 3'b110;
        rom_memory[48305] = 3'b111;
        rom_memory[48306] = 3'b111;
        rom_memory[48307] = 3'b110;
        rom_memory[48308] = 3'b000;
        rom_memory[48309] = 3'b000;
        rom_memory[48310] = 3'b000;
        rom_memory[48311] = 3'b000;
        rom_memory[48312] = 3'b100;
        rom_memory[48313] = 3'b111;
        rom_memory[48314] = 3'b111;
        rom_memory[48315] = 3'b111;
        rom_memory[48316] = 3'b111;
        rom_memory[48317] = 3'b111;
        rom_memory[48318] = 3'b111;
        rom_memory[48319] = 3'b111;
        rom_memory[48320] = 3'b111;
        rom_memory[48321] = 3'b111;
        rom_memory[48322] = 3'b100;
        rom_memory[48323] = 3'b100;
        rom_memory[48324] = 3'b100;
        rom_memory[48325] = 3'b100;
        rom_memory[48326] = 3'b100;
        rom_memory[48327] = 3'b110;
        rom_memory[48328] = 3'b111;
        rom_memory[48329] = 3'b110;
        rom_memory[48330] = 3'b110;
        rom_memory[48331] = 3'b110;
        rom_memory[48332] = 3'b110;
        rom_memory[48333] = 3'b110;
        rom_memory[48334] = 3'b110;
        rom_memory[48335] = 3'b110;
        rom_memory[48336] = 3'b110;
        rom_memory[48337] = 3'b110;
        rom_memory[48338] = 3'b110;
        rom_memory[48339] = 3'b110;
        rom_memory[48340] = 3'b110;
        rom_memory[48341] = 3'b110;
        rom_memory[48342] = 3'b110;
        rom_memory[48343] = 3'b110;
        rom_memory[48344] = 3'b100;
        rom_memory[48345] = 3'b000;
        rom_memory[48346] = 3'b000;
        rom_memory[48347] = 3'b000;
        rom_memory[48348] = 3'b100;
        rom_memory[48349] = 3'b110;
        rom_memory[48350] = 3'b111;
        rom_memory[48351] = 3'b111;
        rom_memory[48352] = 3'b111;
        rom_memory[48353] = 3'b111;
        rom_memory[48354] = 3'b101;
        rom_memory[48355] = 3'b111;
        rom_memory[48356] = 3'b111;
        rom_memory[48357] = 3'b111;
        rom_memory[48358] = 3'b111;
        rom_memory[48359] = 3'b111;
        rom_memory[48360] = 3'b110;
        rom_memory[48361] = 3'b110;
        rom_memory[48362] = 3'b110;
        rom_memory[48363] = 3'b110;
        rom_memory[48364] = 3'b110;
        rom_memory[48365] = 3'b110;
        rom_memory[48366] = 3'b110;
        rom_memory[48367] = 3'b110;
        rom_memory[48368] = 3'b110;
        rom_memory[48369] = 3'b110;
        rom_memory[48370] = 3'b110;
        rom_memory[48371] = 3'b110;
        rom_memory[48372] = 3'b110;
        rom_memory[48373] = 3'b110;
        rom_memory[48374] = 3'b110;
        rom_memory[48375] = 3'b110;
        rom_memory[48376] = 3'b110;
        rom_memory[48377] = 3'b110;
        rom_memory[48378] = 3'b110;
        rom_memory[48379] = 3'b110;
        rom_memory[48380] = 3'b110;
        rom_memory[48381] = 3'b110;
        rom_memory[48382] = 3'b110;
        rom_memory[48383] = 3'b110;
        rom_memory[48384] = 3'b110;
        rom_memory[48385] = 3'b110;
        rom_memory[48386] = 3'b110;
        rom_memory[48387] = 3'b110;
        rom_memory[48388] = 3'b110;
        rom_memory[48389] = 3'b110;
        rom_memory[48390] = 3'b110;
        rom_memory[48391] = 3'b110;
        rom_memory[48392] = 3'b110;
        rom_memory[48393] = 3'b110;
        rom_memory[48394] = 3'b110;
        rom_memory[48395] = 3'b110;
        rom_memory[48396] = 3'b110;
        rom_memory[48397] = 3'b110;
        rom_memory[48398] = 3'b110;
        rom_memory[48399] = 3'b110;
        rom_memory[48400] = 3'b110;
        rom_memory[48401] = 3'b110;
        rom_memory[48402] = 3'b110;
        rom_memory[48403] = 3'b110;
        rom_memory[48404] = 3'b110;
        rom_memory[48405] = 3'b110;
        rom_memory[48406] = 3'b110;
        rom_memory[48407] = 3'b110;
        rom_memory[48408] = 3'b110;
        rom_memory[48409] = 3'b110;
        rom_memory[48410] = 3'b110;
        rom_memory[48411] = 3'b110;
        rom_memory[48412] = 3'b110;
        rom_memory[48413] = 3'b110;
        rom_memory[48414] = 3'b110;
        rom_memory[48415] = 3'b110;
        rom_memory[48416] = 3'b110;
        rom_memory[48417] = 3'b110;
        rom_memory[48418] = 3'b110;
        rom_memory[48419] = 3'b110;
        rom_memory[48420] = 3'b110;
        rom_memory[48421] = 3'b110;
        rom_memory[48422] = 3'b110;
        rom_memory[48423] = 3'b110;
        rom_memory[48424] = 3'b110;
        rom_memory[48425] = 3'b110;
        rom_memory[48426] = 3'b110;
        rom_memory[48427] = 3'b110;
        rom_memory[48428] = 3'b110;
        rom_memory[48429] = 3'b110;
        rom_memory[48430] = 3'b110;
        rom_memory[48431] = 3'b110;
        rom_memory[48432] = 3'b110;
        rom_memory[48433] = 3'b110;
        rom_memory[48434] = 3'b110;
        rom_memory[48435] = 3'b110;
        rom_memory[48436] = 3'b110;
        rom_memory[48437] = 3'b110;
        rom_memory[48438] = 3'b110;
        rom_memory[48439] = 3'b110;
        rom_memory[48440] = 3'b110;
        rom_memory[48441] = 3'b110;
        rom_memory[48442] = 3'b110;
        rom_memory[48443] = 3'b110;
        rom_memory[48444] = 3'b110;
        rom_memory[48445] = 3'b110;
        rom_memory[48446] = 3'b110;
        rom_memory[48447] = 3'b110;
        rom_memory[48448] = 3'b110;
        rom_memory[48449] = 3'b110;
        rom_memory[48450] = 3'b110;
        rom_memory[48451] = 3'b110;
        rom_memory[48452] = 3'b110;
        rom_memory[48453] = 3'b110;
        rom_memory[48454] = 3'b110;
        rom_memory[48455] = 3'b110;
        rom_memory[48456] = 3'b110;
        rom_memory[48457] = 3'b110;
        rom_memory[48458] = 3'b110;
        rom_memory[48459] = 3'b110;
        rom_memory[48460] = 3'b110;
        rom_memory[48461] = 3'b110;
        rom_memory[48462] = 3'b110;
        rom_memory[48463] = 3'b110;
        rom_memory[48464] = 3'b110;
        rom_memory[48465] = 3'b110;
        rom_memory[48466] = 3'b110;
        rom_memory[48467] = 3'b110;
        rom_memory[48468] = 3'b110;
        rom_memory[48469] = 3'b110;
        rom_memory[48470] = 3'b110;
        rom_memory[48471] = 3'b110;
        rom_memory[48472] = 3'b110;
        rom_memory[48473] = 3'b110;
        rom_memory[48474] = 3'b110;
        rom_memory[48475] = 3'b110;
        rom_memory[48476] = 3'b110;
        rom_memory[48477] = 3'b110;
        rom_memory[48478] = 3'b110;
        rom_memory[48479] = 3'b110;
        rom_memory[48480] = 3'b110;
        rom_memory[48481] = 3'b110;
        rom_memory[48482] = 3'b110;
        rom_memory[48483] = 3'b110;
        rom_memory[48484] = 3'b110;
        rom_memory[48485] = 3'b110;
        rom_memory[48486] = 3'b111;
        rom_memory[48487] = 3'b111;
        rom_memory[48488] = 3'b111;
        rom_memory[48489] = 3'b111;
        rom_memory[48490] = 3'b111;
        rom_memory[48491] = 3'b111;
        rom_memory[48492] = 3'b111;
        rom_memory[48493] = 3'b111;
        rom_memory[48494] = 3'b111;
        rom_memory[48495] = 3'b110;
        rom_memory[48496] = 3'b110;
        rom_memory[48497] = 3'b110;
        rom_memory[48498] = 3'b110;
        rom_memory[48499] = 3'b110;
        rom_memory[48500] = 3'b110;
        rom_memory[48501] = 3'b110;
        rom_memory[48502] = 3'b110;
        rom_memory[48503] = 3'b110;
        rom_memory[48504] = 3'b110;
        rom_memory[48505] = 3'b110;
        rom_memory[48506] = 3'b110;
        rom_memory[48507] = 3'b110;
        rom_memory[48508] = 3'b110;
        rom_memory[48509] = 3'b110;
        rom_memory[48510] = 3'b110;
        rom_memory[48511] = 3'b110;
        rom_memory[48512] = 3'b110;
        rom_memory[48513] = 3'b110;
        rom_memory[48514] = 3'b110;
        rom_memory[48515] = 3'b110;
        rom_memory[48516] = 3'b110;
        rom_memory[48517] = 3'b110;
        rom_memory[48518] = 3'b110;
        rom_memory[48519] = 3'b110;
        rom_memory[48520] = 3'b110;
        rom_memory[48521] = 3'b110;
        rom_memory[48522] = 3'b110;
        rom_memory[48523] = 3'b110;
        rom_memory[48524] = 3'b110;
        rom_memory[48525] = 3'b111;
        rom_memory[48526] = 3'b110;
        rom_memory[48527] = 3'b110;
        rom_memory[48528] = 3'b110;
        rom_memory[48529] = 3'b110;
        rom_memory[48530] = 3'b110;
        rom_memory[48531] = 3'b110;
        rom_memory[48532] = 3'b110;
        rom_memory[48533] = 3'b110;
        rom_memory[48534] = 3'b111;
        rom_memory[48535] = 3'b111;
        rom_memory[48536] = 3'b111;
        rom_memory[48537] = 3'b111;
        rom_memory[48538] = 3'b111;
        rom_memory[48539] = 3'b110;
        rom_memory[48540] = 3'b110;
        rom_memory[48541] = 3'b110;
        rom_memory[48542] = 3'b110;
        rom_memory[48543] = 3'b111;
        rom_memory[48544] = 3'b110;
        rom_memory[48545] = 3'b111;
        rom_memory[48546] = 3'b110;
        rom_memory[48547] = 3'b110;
        rom_memory[48548] = 3'b000;
        rom_memory[48549] = 3'b000;
        rom_memory[48550] = 3'b111;
        rom_memory[48551] = 3'b100;
        rom_memory[48552] = 3'b000;
        rom_memory[48553] = 3'b100;
        rom_memory[48554] = 3'b111;
        rom_memory[48555] = 3'b111;
        rom_memory[48556] = 3'b111;
        rom_memory[48557] = 3'b100;
        rom_memory[48558] = 3'b100;
        rom_memory[48559] = 3'b100;
        rom_memory[48560] = 3'b110;
        rom_memory[48561] = 3'b110;
        rom_memory[48562] = 3'b110;
        rom_memory[48563] = 3'b110;
        rom_memory[48564] = 3'b100;
        rom_memory[48565] = 3'b100;
        rom_memory[48566] = 3'b100;
        rom_memory[48567] = 3'b111;
        rom_memory[48568] = 3'b111;
        rom_memory[48569] = 3'b110;
        rom_memory[48570] = 3'b110;
        rom_memory[48571] = 3'b110;
        rom_memory[48572] = 3'b110;
        rom_memory[48573] = 3'b110;
        rom_memory[48574] = 3'b110;
        rom_memory[48575] = 3'b110;
        rom_memory[48576] = 3'b110;
        rom_memory[48577] = 3'b110;
        rom_memory[48578] = 3'b110;
        rom_memory[48579] = 3'b110;
        rom_memory[48580] = 3'b110;
        rom_memory[48581] = 3'b110;
        rom_memory[48582] = 3'b110;
        rom_memory[48583] = 3'b110;
        rom_memory[48584] = 3'b110;
        rom_memory[48585] = 3'b100;
        rom_memory[48586] = 3'b100;
        rom_memory[48587] = 3'b000;
        rom_memory[48588] = 3'b100;
        rom_memory[48589] = 3'b100;
        rom_memory[48590] = 3'b111;
        rom_memory[48591] = 3'b111;
        rom_memory[48592] = 3'b111;
        rom_memory[48593] = 3'b111;
        rom_memory[48594] = 3'b111;
        rom_memory[48595] = 3'b111;
        rom_memory[48596] = 3'b111;
        rom_memory[48597] = 3'b111;
        rom_memory[48598] = 3'b111;
        rom_memory[48599] = 3'b111;
        rom_memory[48600] = 3'b111;
        rom_memory[48601] = 3'b110;
        rom_memory[48602] = 3'b110;
        rom_memory[48603] = 3'b110;
        rom_memory[48604] = 3'b110;
        rom_memory[48605] = 3'b110;
        rom_memory[48606] = 3'b110;
        rom_memory[48607] = 3'b110;
        rom_memory[48608] = 3'b110;
        rom_memory[48609] = 3'b110;
        rom_memory[48610] = 3'b110;
        rom_memory[48611] = 3'b110;
        rom_memory[48612] = 3'b110;
        rom_memory[48613] = 3'b110;
        rom_memory[48614] = 3'b110;
        rom_memory[48615] = 3'b110;
        rom_memory[48616] = 3'b110;
        rom_memory[48617] = 3'b110;
        rom_memory[48618] = 3'b110;
        rom_memory[48619] = 3'b110;
        rom_memory[48620] = 3'b110;
        rom_memory[48621] = 3'b110;
        rom_memory[48622] = 3'b110;
        rom_memory[48623] = 3'b110;
        rom_memory[48624] = 3'b110;
        rom_memory[48625] = 3'b110;
        rom_memory[48626] = 3'b110;
        rom_memory[48627] = 3'b110;
        rom_memory[48628] = 3'b110;
        rom_memory[48629] = 3'b110;
        rom_memory[48630] = 3'b110;
        rom_memory[48631] = 3'b110;
        rom_memory[48632] = 3'b110;
        rom_memory[48633] = 3'b110;
        rom_memory[48634] = 3'b110;
        rom_memory[48635] = 3'b110;
        rom_memory[48636] = 3'b110;
        rom_memory[48637] = 3'b110;
        rom_memory[48638] = 3'b110;
        rom_memory[48639] = 3'b110;
        rom_memory[48640] = 3'b110;
        rom_memory[48641] = 3'b110;
        rom_memory[48642] = 3'b110;
        rom_memory[48643] = 3'b110;
        rom_memory[48644] = 3'b110;
        rom_memory[48645] = 3'b110;
        rom_memory[48646] = 3'b110;
        rom_memory[48647] = 3'b110;
        rom_memory[48648] = 3'b110;
        rom_memory[48649] = 3'b110;
        rom_memory[48650] = 3'b110;
        rom_memory[48651] = 3'b110;
        rom_memory[48652] = 3'b110;
        rom_memory[48653] = 3'b110;
        rom_memory[48654] = 3'b110;
        rom_memory[48655] = 3'b110;
        rom_memory[48656] = 3'b110;
        rom_memory[48657] = 3'b110;
        rom_memory[48658] = 3'b110;
        rom_memory[48659] = 3'b110;
        rom_memory[48660] = 3'b110;
        rom_memory[48661] = 3'b110;
        rom_memory[48662] = 3'b110;
        rom_memory[48663] = 3'b110;
        rom_memory[48664] = 3'b110;
        rom_memory[48665] = 3'b110;
        rom_memory[48666] = 3'b110;
        rom_memory[48667] = 3'b110;
        rom_memory[48668] = 3'b110;
        rom_memory[48669] = 3'b110;
        rom_memory[48670] = 3'b110;
        rom_memory[48671] = 3'b110;
        rom_memory[48672] = 3'b110;
        rom_memory[48673] = 3'b110;
        rom_memory[48674] = 3'b110;
        rom_memory[48675] = 3'b110;
        rom_memory[48676] = 3'b110;
        rom_memory[48677] = 3'b110;
        rom_memory[48678] = 3'b110;
        rom_memory[48679] = 3'b110;
        rom_memory[48680] = 3'b110;
        rom_memory[48681] = 3'b110;
        rom_memory[48682] = 3'b110;
        rom_memory[48683] = 3'b110;
        rom_memory[48684] = 3'b110;
        rom_memory[48685] = 3'b110;
        rom_memory[48686] = 3'b110;
        rom_memory[48687] = 3'b110;
        rom_memory[48688] = 3'b110;
        rom_memory[48689] = 3'b110;
        rom_memory[48690] = 3'b110;
        rom_memory[48691] = 3'b110;
        rom_memory[48692] = 3'b110;
        rom_memory[48693] = 3'b110;
        rom_memory[48694] = 3'b110;
        rom_memory[48695] = 3'b110;
        rom_memory[48696] = 3'b110;
        rom_memory[48697] = 3'b110;
        rom_memory[48698] = 3'b110;
        rom_memory[48699] = 3'b110;
        rom_memory[48700] = 3'b110;
        rom_memory[48701] = 3'b110;
        rom_memory[48702] = 3'b110;
        rom_memory[48703] = 3'b110;
        rom_memory[48704] = 3'b110;
        rom_memory[48705] = 3'b110;
        rom_memory[48706] = 3'b110;
        rom_memory[48707] = 3'b110;
        rom_memory[48708] = 3'b110;
        rom_memory[48709] = 3'b110;
        rom_memory[48710] = 3'b110;
        rom_memory[48711] = 3'b110;
        rom_memory[48712] = 3'b110;
        rom_memory[48713] = 3'b110;
        rom_memory[48714] = 3'b110;
        rom_memory[48715] = 3'b110;
        rom_memory[48716] = 3'b110;
        rom_memory[48717] = 3'b110;
        rom_memory[48718] = 3'b110;
        rom_memory[48719] = 3'b110;
        rom_memory[48720] = 3'b110;
        rom_memory[48721] = 3'b110;
        rom_memory[48722] = 3'b110;
        rom_memory[48723] = 3'b110;
        rom_memory[48724] = 3'b110;
        rom_memory[48725] = 3'b110;
        rom_memory[48726] = 3'b110;
        rom_memory[48727] = 3'b111;
        rom_memory[48728] = 3'b111;
        rom_memory[48729] = 3'b111;
        rom_memory[48730] = 3'b111;
        rom_memory[48731] = 3'b111;
        rom_memory[48732] = 3'b111;
        rom_memory[48733] = 3'b111;
        rom_memory[48734] = 3'b110;
        rom_memory[48735] = 3'b110;
        rom_memory[48736] = 3'b110;
        rom_memory[48737] = 3'b110;
        rom_memory[48738] = 3'b110;
        rom_memory[48739] = 3'b110;
        rom_memory[48740] = 3'b110;
        rom_memory[48741] = 3'b110;
        rom_memory[48742] = 3'b110;
        rom_memory[48743] = 3'b110;
        rom_memory[48744] = 3'b110;
        rom_memory[48745] = 3'b110;
        rom_memory[48746] = 3'b110;
        rom_memory[48747] = 3'b110;
        rom_memory[48748] = 3'b110;
        rom_memory[48749] = 3'b110;
        rom_memory[48750] = 3'b110;
        rom_memory[48751] = 3'b110;
        rom_memory[48752] = 3'b110;
        rom_memory[48753] = 3'b110;
        rom_memory[48754] = 3'b110;
        rom_memory[48755] = 3'b110;
        rom_memory[48756] = 3'b110;
        rom_memory[48757] = 3'b110;
        rom_memory[48758] = 3'b110;
        rom_memory[48759] = 3'b110;
        rom_memory[48760] = 3'b110;
        rom_memory[48761] = 3'b110;
        rom_memory[48762] = 3'b110;
        rom_memory[48763] = 3'b110;
        rom_memory[48764] = 3'b110;
        rom_memory[48765] = 3'b111;
        rom_memory[48766] = 3'b110;
        rom_memory[48767] = 3'b110;
        rom_memory[48768] = 3'b110;
        rom_memory[48769] = 3'b110;
        rom_memory[48770] = 3'b110;
        rom_memory[48771] = 3'b010;
        rom_memory[48772] = 3'b110;
        rom_memory[48773] = 3'b110;
        rom_memory[48774] = 3'b111;
        rom_memory[48775] = 3'b111;
        rom_memory[48776] = 3'b111;
        rom_memory[48777] = 3'b111;
        rom_memory[48778] = 3'b110;
        rom_memory[48779] = 3'b110;
        rom_memory[48780] = 3'b110;
        rom_memory[48781] = 3'b110;
        rom_memory[48782] = 3'b111;
        rom_memory[48783] = 3'b111;
        rom_memory[48784] = 3'b110;
        rom_memory[48785] = 3'b111;
        rom_memory[48786] = 3'b111;
        rom_memory[48787] = 3'b110;
        rom_memory[48788] = 3'b000;
        rom_memory[48789] = 3'b000;
        rom_memory[48790] = 3'b100;
        rom_memory[48791] = 3'b111;
        rom_memory[48792] = 3'b000;
        rom_memory[48793] = 3'b111;
        rom_memory[48794] = 3'b111;
        rom_memory[48795] = 3'b111;
        rom_memory[48796] = 3'b100;
        rom_memory[48797] = 3'b100;
        rom_memory[48798] = 3'b100;
        rom_memory[48799] = 3'b100;
        rom_memory[48800] = 3'b100;
        rom_memory[48801] = 3'b100;
        rom_memory[48802] = 3'b100;
        rom_memory[48803] = 3'b100;
        rom_memory[48804] = 3'b100;
        rom_memory[48805] = 3'b100;
        rom_memory[48806] = 3'b110;
        rom_memory[48807] = 3'b111;
        rom_memory[48808] = 3'b111;
        rom_memory[48809] = 3'b110;
        rom_memory[48810] = 3'b110;
        rom_memory[48811] = 3'b110;
        rom_memory[48812] = 3'b110;
        rom_memory[48813] = 3'b110;
        rom_memory[48814] = 3'b110;
        rom_memory[48815] = 3'b110;
        rom_memory[48816] = 3'b110;
        rom_memory[48817] = 3'b110;
        rom_memory[48818] = 3'b110;
        rom_memory[48819] = 3'b110;
        rom_memory[48820] = 3'b110;
        rom_memory[48821] = 3'b110;
        rom_memory[48822] = 3'b110;
        rom_memory[48823] = 3'b110;
        rom_memory[48824] = 3'b110;
        rom_memory[48825] = 3'b110;
        rom_memory[48826] = 3'b100;
        rom_memory[48827] = 3'b100;
        rom_memory[48828] = 3'b100;
        rom_memory[48829] = 3'b100;
        rom_memory[48830] = 3'b111;
        rom_memory[48831] = 3'b111;
        rom_memory[48832] = 3'b111;
        rom_memory[48833] = 3'b111;
        rom_memory[48834] = 3'b111;
        rom_memory[48835] = 3'b111;
        rom_memory[48836] = 3'b111;
        rom_memory[48837] = 3'b111;
        rom_memory[48838] = 3'b111;
        rom_memory[48839] = 3'b111;
        rom_memory[48840] = 3'b111;
        rom_memory[48841] = 3'b110;
        rom_memory[48842] = 3'b110;
        rom_memory[48843] = 3'b110;
        rom_memory[48844] = 3'b110;
        rom_memory[48845] = 3'b110;
        rom_memory[48846] = 3'b110;
        rom_memory[48847] = 3'b110;
        rom_memory[48848] = 3'b110;
        rom_memory[48849] = 3'b110;
        rom_memory[48850] = 3'b110;
        rom_memory[48851] = 3'b110;
        rom_memory[48852] = 3'b110;
        rom_memory[48853] = 3'b110;
        rom_memory[48854] = 3'b110;
        rom_memory[48855] = 3'b110;
        rom_memory[48856] = 3'b110;
        rom_memory[48857] = 3'b110;
        rom_memory[48858] = 3'b110;
        rom_memory[48859] = 3'b110;
        rom_memory[48860] = 3'b110;
        rom_memory[48861] = 3'b110;
        rom_memory[48862] = 3'b110;
        rom_memory[48863] = 3'b110;
        rom_memory[48864] = 3'b110;
        rom_memory[48865] = 3'b110;
        rom_memory[48866] = 3'b110;
        rom_memory[48867] = 3'b110;
        rom_memory[48868] = 3'b110;
        rom_memory[48869] = 3'b110;
        rom_memory[48870] = 3'b110;
        rom_memory[48871] = 3'b110;
        rom_memory[48872] = 3'b110;
        rom_memory[48873] = 3'b110;
        rom_memory[48874] = 3'b110;
        rom_memory[48875] = 3'b110;
        rom_memory[48876] = 3'b110;
        rom_memory[48877] = 3'b110;
        rom_memory[48878] = 3'b110;
        rom_memory[48879] = 3'b110;
        rom_memory[48880] = 3'b110;
        rom_memory[48881] = 3'b110;
        rom_memory[48882] = 3'b110;
        rom_memory[48883] = 3'b110;
        rom_memory[48884] = 3'b110;
        rom_memory[48885] = 3'b110;
        rom_memory[48886] = 3'b110;
        rom_memory[48887] = 3'b110;
        rom_memory[48888] = 3'b110;
        rom_memory[48889] = 3'b110;
        rom_memory[48890] = 3'b110;
        rom_memory[48891] = 3'b110;
        rom_memory[48892] = 3'b110;
        rom_memory[48893] = 3'b110;
        rom_memory[48894] = 3'b110;
        rom_memory[48895] = 3'b110;
        rom_memory[48896] = 3'b110;
        rom_memory[48897] = 3'b110;
        rom_memory[48898] = 3'b110;
        rom_memory[48899] = 3'b110;
        rom_memory[48900] = 3'b110;
        rom_memory[48901] = 3'b110;
        rom_memory[48902] = 3'b110;
        rom_memory[48903] = 3'b110;
        rom_memory[48904] = 3'b110;
        rom_memory[48905] = 3'b110;
        rom_memory[48906] = 3'b110;
        rom_memory[48907] = 3'b110;
        rom_memory[48908] = 3'b110;
        rom_memory[48909] = 3'b110;
        rom_memory[48910] = 3'b110;
        rom_memory[48911] = 3'b110;
        rom_memory[48912] = 3'b110;
        rom_memory[48913] = 3'b110;
        rom_memory[48914] = 3'b110;
        rom_memory[48915] = 3'b110;
        rom_memory[48916] = 3'b110;
        rom_memory[48917] = 3'b110;
        rom_memory[48918] = 3'b110;
        rom_memory[48919] = 3'b110;
        rom_memory[48920] = 3'b110;
        rom_memory[48921] = 3'b110;
        rom_memory[48922] = 3'b110;
        rom_memory[48923] = 3'b110;
        rom_memory[48924] = 3'b110;
        rom_memory[48925] = 3'b110;
        rom_memory[48926] = 3'b110;
        rom_memory[48927] = 3'b110;
        rom_memory[48928] = 3'b110;
        rom_memory[48929] = 3'b110;
        rom_memory[48930] = 3'b110;
        rom_memory[48931] = 3'b110;
        rom_memory[48932] = 3'b110;
        rom_memory[48933] = 3'b110;
        rom_memory[48934] = 3'b110;
        rom_memory[48935] = 3'b110;
        rom_memory[48936] = 3'b110;
        rom_memory[48937] = 3'b110;
        rom_memory[48938] = 3'b110;
        rom_memory[48939] = 3'b110;
        rom_memory[48940] = 3'b110;
        rom_memory[48941] = 3'b110;
        rom_memory[48942] = 3'b110;
        rom_memory[48943] = 3'b110;
        rom_memory[48944] = 3'b110;
        rom_memory[48945] = 3'b110;
        rom_memory[48946] = 3'b110;
        rom_memory[48947] = 3'b110;
        rom_memory[48948] = 3'b110;
        rom_memory[48949] = 3'b110;
        rom_memory[48950] = 3'b110;
        rom_memory[48951] = 3'b110;
        rom_memory[48952] = 3'b110;
        rom_memory[48953] = 3'b110;
        rom_memory[48954] = 3'b110;
        rom_memory[48955] = 3'b110;
        rom_memory[48956] = 3'b110;
        rom_memory[48957] = 3'b110;
        rom_memory[48958] = 3'b110;
        rom_memory[48959] = 3'b110;
        rom_memory[48960] = 3'b110;
        rom_memory[48961] = 3'b110;
        rom_memory[48962] = 3'b110;
        rom_memory[48963] = 3'b110;
        rom_memory[48964] = 3'b110;
        rom_memory[48965] = 3'b110;
        rom_memory[48966] = 3'b110;
        rom_memory[48967] = 3'b110;
        rom_memory[48968] = 3'b111;
        rom_memory[48969] = 3'b111;
        rom_memory[48970] = 3'b111;
        rom_memory[48971] = 3'b111;
        rom_memory[48972] = 3'b111;
        rom_memory[48973] = 3'b111;
        rom_memory[48974] = 3'b110;
        rom_memory[48975] = 3'b110;
        rom_memory[48976] = 3'b110;
        rom_memory[48977] = 3'b110;
        rom_memory[48978] = 3'b110;
        rom_memory[48979] = 3'b110;
        rom_memory[48980] = 3'b110;
        rom_memory[48981] = 3'b110;
        rom_memory[48982] = 3'b110;
        rom_memory[48983] = 3'b110;
        rom_memory[48984] = 3'b110;
        rom_memory[48985] = 3'b110;
        rom_memory[48986] = 3'b110;
        rom_memory[48987] = 3'b110;
        rom_memory[48988] = 3'b110;
        rom_memory[48989] = 3'b110;
        rom_memory[48990] = 3'b110;
        rom_memory[48991] = 3'b110;
        rom_memory[48992] = 3'b110;
        rom_memory[48993] = 3'b110;
        rom_memory[48994] = 3'b110;
        rom_memory[48995] = 3'b110;
        rom_memory[48996] = 3'b110;
        rom_memory[48997] = 3'b110;
        rom_memory[48998] = 3'b110;
        rom_memory[48999] = 3'b110;
        rom_memory[49000] = 3'b110;
        rom_memory[49001] = 3'b110;
        rom_memory[49002] = 3'b110;
        rom_memory[49003] = 3'b110;
        rom_memory[49004] = 3'b110;
        rom_memory[49005] = 3'b111;
        rom_memory[49006] = 3'b111;
        rom_memory[49007] = 3'b110;
        rom_memory[49008] = 3'b110;
        rom_memory[49009] = 3'b110;
        rom_memory[49010] = 3'b110;
        rom_memory[49011] = 3'b110;
        rom_memory[49012] = 3'b110;
        rom_memory[49013] = 3'b110;
        rom_memory[49014] = 3'b111;
        rom_memory[49015] = 3'b110;
        rom_memory[49016] = 3'b111;
        rom_memory[49017] = 3'b111;
        rom_memory[49018] = 3'b110;
        rom_memory[49019] = 3'b110;
        rom_memory[49020] = 3'b110;
        rom_memory[49021] = 3'b110;
        rom_memory[49022] = 3'b111;
        rom_memory[49023] = 3'b111;
        rom_memory[49024] = 3'b110;
        rom_memory[49025] = 3'b111;
        rom_memory[49026] = 3'b111;
        rom_memory[49027] = 3'b111;
        rom_memory[49028] = 3'b100;
        rom_memory[49029] = 3'b100;
        rom_memory[49030] = 3'b111;
        rom_memory[49031] = 3'b111;
        rom_memory[49032] = 3'b111;
        rom_memory[49033] = 3'b111;
        rom_memory[49034] = 3'b111;
        rom_memory[49035] = 3'b100;
        rom_memory[49036] = 3'b100;
        rom_memory[49037] = 3'b000;
        rom_memory[49038] = 3'b000;
        rom_memory[49039] = 3'b000;
        rom_memory[49040] = 3'b100;
        rom_memory[49041] = 3'b100;
        rom_memory[49042] = 3'b100;
        rom_memory[49043] = 3'b100;
        rom_memory[49044] = 3'b100;
        rom_memory[49045] = 3'b100;
        rom_memory[49046] = 3'b111;
        rom_memory[49047] = 3'b111;
        rom_memory[49048] = 3'b111;
        rom_memory[49049] = 3'b110;
        rom_memory[49050] = 3'b110;
        rom_memory[49051] = 3'b100;
        rom_memory[49052] = 3'b110;
        rom_memory[49053] = 3'b110;
        rom_memory[49054] = 3'b110;
        rom_memory[49055] = 3'b110;
        rom_memory[49056] = 3'b110;
        rom_memory[49057] = 3'b110;
        rom_memory[49058] = 3'b110;
        rom_memory[49059] = 3'b110;
        rom_memory[49060] = 3'b110;
        rom_memory[49061] = 3'b110;
        rom_memory[49062] = 3'b110;
        rom_memory[49063] = 3'b110;
        rom_memory[49064] = 3'b110;
        rom_memory[49065] = 3'b110;
        rom_memory[49066] = 3'b110;
        rom_memory[49067] = 3'b100;
        rom_memory[49068] = 3'b100;
        rom_memory[49069] = 3'b100;
        rom_memory[49070] = 3'b100;
        rom_memory[49071] = 3'b100;
        rom_memory[49072] = 3'b101;
        rom_memory[49073] = 3'b111;
        rom_memory[49074] = 3'b111;
        rom_memory[49075] = 3'b111;
        rom_memory[49076] = 3'b111;
        rom_memory[49077] = 3'b111;
        rom_memory[49078] = 3'b111;
        rom_memory[49079] = 3'b111;
        rom_memory[49080] = 3'b111;
        rom_memory[49081] = 3'b110;
        rom_memory[49082] = 3'b110;
        rom_memory[49083] = 3'b110;
        rom_memory[49084] = 3'b110;
        rom_memory[49085] = 3'b110;
        rom_memory[49086] = 3'b110;
        rom_memory[49087] = 3'b110;
        rom_memory[49088] = 3'b110;
        rom_memory[49089] = 3'b110;
        rom_memory[49090] = 3'b110;
        rom_memory[49091] = 3'b110;
        rom_memory[49092] = 3'b110;
        rom_memory[49093] = 3'b110;
        rom_memory[49094] = 3'b110;
        rom_memory[49095] = 3'b110;
        rom_memory[49096] = 3'b110;
        rom_memory[49097] = 3'b110;
        rom_memory[49098] = 3'b110;
        rom_memory[49099] = 3'b110;
        rom_memory[49100] = 3'b110;
        rom_memory[49101] = 3'b110;
        rom_memory[49102] = 3'b110;
        rom_memory[49103] = 3'b110;
        rom_memory[49104] = 3'b110;
        rom_memory[49105] = 3'b110;
        rom_memory[49106] = 3'b110;
        rom_memory[49107] = 3'b110;
        rom_memory[49108] = 3'b110;
        rom_memory[49109] = 3'b110;
        rom_memory[49110] = 3'b110;
        rom_memory[49111] = 3'b110;
        rom_memory[49112] = 3'b110;
        rom_memory[49113] = 3'b110;
        rom_memory[49114] = 3'b110;
        rom_memory[49115] = 3'b110;
        rom_memory[49116] = 3'b110;
        rom_memory[49117] = 3'b110;
        rom_memory[49118] = 3'b110;
        rom_memory[49119] = 3'b110;
        rom_memory[49120] = 3'b110;
        rom_memory[49121] = 3'b110;
        rom_memory[49122] = 3'b110;
        rom_memory[49123] = 3'b110;
        rom_memory[49124] = 3'b110;
        rom_memory[49125] = 3'b110;
        rom_memory[49126] = 3'b110;
        rom_memory[49127] = 3'b110;
        rom_memory[49128] = 3'b110;
        rom_memory[49129] = 3'b110;
        rom_memory[49130] = 3'b110;
        rom_memory[49131] = 3'b110;
        rom_memory[49132] = 3'b110;
        rom_memory[49133] = 3'b110;
        rom_memory[49134] = 3'b110;
        rom_memory[49135] = 3'b110;
        rom_memory[49136] = 3'b110;
        rom_memory[49137] = 3'b110;
        rom_memory[49138] = 3'b110;
        rom_memory[49139] = 3'b110;
        rom_memory[49140] = 3'b110;
        rom_memory[49141] = 3'b110;
        rom_memory[49142] = 3'b110;
        rom_memory[49143] = 3'b110;
        rom_memory[49144] = 3'b110;
        rom_memory[49145] = 3'b110;
        rom_memory[49146] = 3'b110;
        rom_memory[49147] = 3'b110;
        rom_memory[49148] = 3'b110;
        rom_memory[49149] = 3'b110;
        rom_memory[49150] = 3'b110;
        rom_memory[49151] = 3'b110;
        rom_memory[49152] = 3'b110;
        rom_memory[49153] = 3'b110;
        rom_memory[49154] = 3'b110;
        rom_memory[49155] = 3'b110;
        rom_memory[49156] = 3'b110;
        rom_memory[49157] = 3'b110;
        rom_memory[49158] = 3'b110;
        rom_memory[49159] = 3'b110;
        rom_memory[49160] = 3'b110;
        rom_memory[49161] = 3'b110;
        rom_memory[49162] = 3'b110;
        rom_memory[49163] = 3'b110;
        rom_memory[49164] = 3'b110;
        rom_memory[49165] = 3'b110;
        rom_memory[49166] = 3'b110;
        rom_memory[49167] = 3'b110;
        rom_memory[49168] = 3'b110;
        rom_memory[49169] = 3'b110;
        rom_memory[49170] = 3'b110;
        rom_memory[49171] = 3'b110;
        rom_memory[49172] = 3'b110;
        rom_memory[49173] = 3'b110;
        rom_memory[49174] = 3'b110;
        rom_memory[49175] = 3'b110;
        rom_memory[49176] = 3'b110;
        rom_memory[49177] = 3'b110;
        rom_memory[49178] = 3'b110;
        rom_memory[49179] = 3'b110;
        rom_memory[49180] = 3'b110;
        rom_memory[49181] = 3'b110;
        rom_memory[49182] = 3'b110;
        rom_memory[49183] = 3'b110;
        rom_memory[49184] = 3'b110;
        rom_memory[49185] = 3'b110;
        rom_memory[49186] = 3'b110;
        rom_memory[49187] = 3'b110;
        rom_memory[49188] = 3'b110;
        rom_memory[49189] = 3'b110;
        rom_memory[49190] = 3'b110;
        rom_memory[49191] = 3'b110;
        rom_memory[49192] = 3'b110;
        rom_memory[49193] = 3'b110;
        rom_memory[49194] = 3'b110;
        rom_memory[49195] = 3'b110;
        rom_memory[49196] = 3'b110;
        rom_memory[49197] = 3'b110;
        rom_memory[49198] = 3'b110;
        rom_memory[49199] = 3'b110;
        rom_memory[49200] = 3'b110;
        rom_memory[49201] = 3'b110;
        rom_memory[49202] = 3'b110;
        rom_memory[49203] = 3'b110;
        rom_memory[49204] = 3'b110;
        rom_memory[49205] = 3'b110;
        rom_memory[49206] = 3'b110;
        rom_memory[49207] = 3'b110;
        rom_memory[49208] = 3'b110;
        rom_memory[49209] = 3'b110;
        rom_memory[49210] = 3'b111;
        rom_memory[49211] = 3'b111;
        rom_memory[49212] = 3'b111;
        rom_memory[49213] = 3'b111;
        rom_memory[49214] = 3'b110;
        rom_memory[49215] = 3'b110;
        rom_memory[49216] = 3'b110;
        rom_memory[49217] = 3'b110;
        rom_memory[49218] = 3'b110;
        rom_memory[49219] = 3'b110;
        rom_memory[49220] = 3'b110;
        rom_memory[49221] = 3'b110;
        rom_memory[49222] = 3'b110;
        rom_memory[49223] = 3'b110;
        rom_memory[49224] = 3'b110;
        rom_memory[49225] = 3'b110;
        rom_memory[49226] = 3'b110;
        rom_memory[49227] = 3'b110;
        rom_memory[49228] = 3'b110;
        rom_memory[49229] = 3'b110;
        rom_memory[49230] = 3'b110;
        rom_memory[49231] = 3'b110;
        rom_memory[49232] = 3'b110;
        rom_memory[49233] = 3'b110;
        rom_memory[49234] = 3'b110;
        rom_memory[49235] = 3'b110;
        rom_memory[49236] = 3'b110;
        rom_memory[49237] = 3'b110;
        rom_memory[49238] = 3'b110;
        rom_memory[49239] = 3'b110;
        rom_memory[49240] = 3'b110;
        rom_memory[49241] = 3'b110;
        rom_memory[49242] = 3'b110;
        rom_memory[49243] = 3'b110;
        rom_memory[49244] = 3'b110;
        rom_memory[49245] = 3'b110;
        rom_memory[49246] = 3'b111;
        rom_memory[49247] = 3'b111;
        rom_memory[49248] = 3'b110;
        rom_memory[49249] = 3'b110;
        rom_memory[49250] = 3'b110;
        rom_memory[49251] = 3'b110;
        rom_memory[49252] = 3'b110;
        rom_memory[49253] = 3'b110;
        rom_memory[49254] = 3'b110;
        rom_memory[49255] = 3'b110;
        rom_memory[49256] = 3'b110;
        rom_memory[49257] = 3'b110;
        rom_memory[49258] = 3'b110;
        rom_memory[49259] = 3'b110;
        rom_memory[49260] = 3'b110;
        rom_memory[49261] = 3'b110;
        rom_memory[49262] = 3'b111;
        rom_memory[49263] = 3'b111;
        rom_memory[49264] = 3'b111;
        rom_memory[49265] = 3'b111;
        rom_memory[49266] = 3'b111;
        rom_memory[49267] = 3'b111;
        rom_memory[49268] = 3'b000;
        rom_memory[49269] = 3'b111;
        rom_memory[49270] = 3'b111;
        rom_memory[49271] = 3'b111;
        rom_memory[49272] = 3'b100;
        rom_memory[49273] = 3'b100;
        rom_memory[49274] = 3'b000;
        rom_memory[49275] = 3'b000;
        rom_memory[49276] = 3'b000;
        rom_memory[49277] = 3'b000;
        rom_memory[49278] = 3'b000;
        rom_memory[49279] = 3'b000;
        rom_memory[49280] = 3'b000;
        rom_memory[49281] = 3'b100;
        rom_memory[49282] = 3'b100;
        rom_memory[49283] = 3'b100;
        rom_memory[49284] = 3'b100;
        rom_memory[49285] = 3'b100;
        rom_memory[49286] = 3'b111;
        rom_memory[49287] = 3'b111;
        rom_memory[49288] = 3'b110;
        rom_memory[49289] = 3'b111;
        rom_memory[49290] = 3'b110;
        rom_memory[49291] = 3'b100;
        rom_memory[49292] = 3'b110;
        rom_memory[49293] = 3'b110;
        rom_memory[49294] = 3'b110;
        rom_memory[49295] = 3'b110;
        rom_memory[49296] = 3'b110;
        rom_memory[49297] = 3'b110;
        rom_memory[49298] = 3'b110;
        rom_memory[49299] = 3'b110;
        rom_memory[49300] = 3'b110;
        rom_memory[49301] = 3'b110;
        rom_memory[49302] = 3'b110;
        rom_memory[49303] = 3'b110;
        rom_memory[49304] = 3'b110;
        rom_memory[49305] = 3'b110;
        rom_memory[49306] = 3'b111;
        rom_memory[49307] = 3'b110;
        rom_memory[49308] = 3'b100;
        rom_memory[49309] = 3'b100;
        rom_memory[49310] = 3'b100;
        rom_memory[49311] = 3'b100;
        rom_memory[49312] = 3'b100;
        rom_memory[49313] = 3'b111;
        rom_memory[49314] = 3'b111;
        rom_memory[49315] = 3'b111;
        rom_memory[49316] = 3'b111;
        rom_memory[49317] = 3'b111;
        rom_memory[49318] = 3'b111;
        rom_memory[49319] = 3'b111;
        rom_memory[49320] = 3'b111;
        rom_memory[49321] = 3'b111;
        rom_memory[49322] = 3'b110;
        rom_memory[49323] = 3'b110;
        rom_memory[49324] = 3'b110;
        rom_memory[49325] = 3'b110;
        rom_memory[49326] = 3'b110;
        rom_memory[49327] = 3'b110;
        rom_memory[49328] = 3'b110;
        rom_memory[49329] = 3'b110;
        rom_memory[49330] = 3'b110;
        rom_memory[49331] = 3'b110;
        rom_memory[49332] = 3'b110;
        rom_memory[49333] = 3'b110;
        rom_memory[49334] = 3'b110;
        rom_memory[49335] = 3'b110;
        rom_memory[49336] = 3'b110;
        rom_memory[49337] = 3'b110;
        rom_memory[49338] = 3'b110;
        rom_memory[49339] = 3'b110;
        rom_memory[49340] = 3'b110;
        rom_memory[49341] = 3'b110;
        rom_memory[49342] = 3'b110;
        rom_memory[49343] = 3'b110;
        rom_memory[49344] = 3'b110;
        rom_memory[49345] = 3'b110;
        rom_memory[49346] = 3'b110;
        rom_memory[49347] = 3'b110;
        rom_memory[49348] = 3'b110;
        rom_memory[49349] = 3'b110;
        rom_memory[49350] = 3'b110;
        rom_memory[49351] = 3'b110;
        rom_memory[49352] = 3'b110;
        rom_memory[49353] = 3'b110;
        rom_memory[49354] = 3'b110;
        rom_memory[49355] = 3'b110;
        rom_memory[49356] = 3'b110;
        rom_memory[49357] = 3'b110;
        rom_memory[49358] = 3'b110;
        rom_memory[49359] = 3'b110;
        rom_memory[49360] = 3'b110;
        rom_memory[49361] = 3'b110;
        rom_memory[49362] = 3'b110;
        rom_memory[49363] = 3'b110;
        rom_memory[49364] = 3'b110;
        rom_memory[49365] = 3'b110;
        rom_memory[49366] = 3'b110;
        rom_memory[49367] = 3'b110;
        rom_memory[49368] = 3'b110;
        rom_memory[49369] = 3'b110;
        rom_memory[49370] = 3'b110;
        rom_memory[49371] = 3'b110;
        rom_memory[49372] = 3'b110;
        rom_memory[49373] = 3'b110;
        rom_memory[49374] = 3'b110;
        rom_memory[49375] = 3'b110;
        rom_memory[49376] = 3'b110;
        rom_memory[49377] = 3'b110;
        rom_memory[49378] = 3'b110;
        rom_memory[49379] = 3'b110;
        rom_memory[49380] = 3'b110;
        rom_memory[49381] = 3'b110;
        rom_memory[49382] = 3'b110;
        rom_memory[49383] = 3'b110;
        rom_memory[49384] = 3'b110;
        rom_memory[49385] = 3'b110;
        rom_memory[49386] = 3'b110;
        rom_memory[49387] = 3'b110;
        rom_memory[49388] = 3'b110;
        rom_memory[49389] = 3'b110;
        rom_memory[49390] = 3'b110;
        rom_memory[49391] = 3'b110;
        rom_memory[49392] = 3'b110;
        rom_memory[49393] = 3'b110;
        rom_memory[49394] = 3'b110;
        rom_memory[49395] = 3'b110;
        rom_memory[49396] = 3'b110;
        rom_memory[49397] = 3'b110;
        rom_memory[49398] = 3'b110;
        rom_memory[49399] = 3'b110;
        rom_memory[49400] = 3'b110;
        rom_memory[49401] = 3'b110;
        rom_memory[49402] = 3'b110;
        rom_memory[49403] = 3'b110;
        rom_memory[49404] = 3'b110;
        rom_memory[49405] = 3'b110;
        rom_memory[49406] = 3'b110;
        rom_memory[49407] = 3'b110;
        rom_memory[49408] = 3'b110;
        rom_memory[49409] = 3'b110;
        rom_memory[49410] = 3'b110;
        rom_memory[49411] = 3'b110;
        rom_memory[49412] = 3'b110;
        rom_memory[49413] = 3'b110;
        rom_memory[49414] = 3'b110;
        rom_memory[49415] = 3'b110;
        rom_memory[49416] = 3'b110;
        rom_memory[49417] = 3'b110;
        rom_memory[49418] = 3'b110;
        rom_memory[49419] = 3'b110;
        rom_memory[49420] = 3'b110;
        rom_memory[49421] = 3'b110;
        rom_memory[49422] = 3'b110;
        rom_memory[49423] = 3'b110;
        rom_memory[49424] = 3'b110;
        rom_memory[49425] = 3'b110;
        rom_memory[49426] = 3'b110;
        rom_memory[49427] = 3'b110;
        rom_memory[49428] = 3'b110;
        rom_memory[49429] = 3'b110;
        rom_memory[49430] = 3'b110;
        rom_memory[49431] = 3'b110;
        rom_memory[49432] = 3'b110;
        rom_memory[49433] = 3'b110;
        rom_memory[49434] = 3'b110;
        rom_memory[49435] = 3'b110;
        rom_memory[49436] = 3'b110;
        rom_memory[49437] = 3'b110;
        rom_memory[49438] = 3'b110;
        rom_memory[49439] = 3'b110;
        rom_memory[49440] = 3'b110;
        rom_memory[49441] = 3'b110;
        rom_memory[49442] = 3'b110;
        rom_memory[49443] = 3'b110;
        rom_memory[49444] = 3'b110;
        rom_memory[49445] = 3'b110;
        rom_memory[49446] = 3'b110;
        rom_memory[49447] = 3'b110;
        rom_memory[49448] = 3'b110;
        rom_memory[49449] = 3'b110;
        rom_memory[49450] = 3'b110;
        rom_memory[49451] = 3'b111;
        rom_memory[49452] = 3'b110;
        rom_memory[49453] = 3'b110;
        rom_memory[49454] = 3'b110;
        rom_memory[49455] = 3'b110;
        rom_memory[49456] = 3'b110;
        rom_memory[49457] = 3'b110;
        rom_memory[49458] = 3'b110;
        rom_memory[49459] = 3'b110;
        rom_memory[49460] = 3'b110;
        rom_memory[49461] = 3'b110;
        rom_memory[49462] = 3'b110;
        rom_memory[49463] = 3'b110;
        rom_memory[49464] = 3'b110;
        rom_memory[49465] = 3'b110;
        rom_memory[49466] = 3'b110;
        rom_memory[49467] = 3'b110;
        rom_memory[49468] = 3'b110;
        rom_memory[49469] = 3'b110;
        rom_memory[49470] = 3'b110;
        rom_memory[49471] = 3'b110;
        rom_memory[49472] = 3'b110;
        rom_memory[49473] = 3'b110;
        rom_memory[49474] = 3'b110;
        rom_memory[49475] = 3'b110;
        rom_memory[49476] = 3'b110;
        rom_memory[49477] = 3'b110;
        rom_memory[49478] = 3'b110;
        rom_memory[49479] = 3'b110;
        rom_memory[49480] = 3'b110;
        rom_memory[49481] = 3'b110;
        rom_memory[49482] = 3'b110;
        rom_memory[49483] = 3'b110;
        rom_memory[49484] = 3'b110;
        rom_memory[49485] = 3'b110;
        rom_memory[49486] = 3'b111;
        rom_memory[49487] = 3'b111;
        rom_memory[49488] = 3'b111;
        rom_memory[49489] = 3'b110;
        rom_memory[49490] = 3'b110;
        rom_memory[49491] = 3'b110;
        rom_memory[49492] = 3'b110;
        rom_memory[49493] = 3'b110;
        rom_memory[49494] = 3'b110;
        rom_memory[49495] = 3'b110;
        rom_memory[49496] = 3'b110;
        rom_memory[49497] = 3'b110;
        rom_memory[49498] = 3'b110;
        rom_memory[49499] = 3'b110;
        rom_memory[49500] = 3'b110;
        rom_memory[49501] = 3'b111;
        rom_memory[49502] = 3'b111;
        rom_memory[49503] = 3'b111;
        rom_memory[49504] = 3'b111;
        rom_memory[49505] = 3'b111;
        rom_memory[49506] = 3'b111;
        rom_memory[49507] = 3'b111;
        rom_memory[49508] = 3'b000;
        rom_memory[49509] = 3'b111;
        rom_memory[49510] = 3'b100;
        rom_memory[49511] = 3'b111;
        rom_memory[49512] = 3'b000;
        rom_memory[49513] = 3'b100;
        rom_memory[49514] = 3'b000;
        rom_memory[49515] = 3'b000;
        rom_memory[49516] = 3'b000;
        rom_memory[49517] = 3'b000;
        rom_memory[49518] = 3'b000;
        rom_memory[49519] = 3'b000;
        rom_memory[49520] = 3'b000;
        rom_memory[49521] = 3'b000;
        rom_memory[49522] = 3'b000;
        rom_memory[49523] = 3'b100;
        rom_memory[49524] = 3'b100;
        rom_memory[49525] = 3'b110;
        rom_memory[49526] = 3'b111;
        rom_memory[49527] = 3'b111;
        rom_memory[49528] = 3'b110;
        rom_memory[49529] = 3'b111;
        rom_memory[49530] = 3'b110;
        rom_memory[49531] = 3'b100;
        rom_memory[49532] = 3'b100;
        rom_memory[49533] = 3'b110;
        rom_memory[49534] = 3'b110;
        rom_memory[49535] = 3'b110;
        rom_memory[49536] = 3'b110;
        rom_memory[49537] = 3'b110;
        rom_memory[49538] = 3'b110;
        rom_memory[49539] = 3'b110;
        rom_memory[49540] = 3'b110;
        rom_memory[49541] = 3'b110;
        rom_memory[49542] = 3'b110;
        rom_memory[49543] = 3'b110;
        rom_memory[49544] = 3'b110;
        rom_memory[49545] = 3'b111;
        rom_memory[49546] = 3'b111;
        rom_memory[49547] = 3'b110;
        rom_memory[49548] = 3'b100;
        rom_memory[49549] = 3'b100;
        rom_memory[49550] = 3'b000;
        rom_memory[49551] = 3'b100;
        rom_memory[49552] = 3'b100;
        rom_memory[49553] = 3'b100;
        rom_memory[49554] = 3'b111;
        rom_memory[49555] = 3'b111;
        rom_memory[49556] = 3'b111;
        rom_memory[49557] = 3'b111;
        rom_memory[49558] = 3'b111;
        rom_memory[49559] = 3'b111;
        rom_memory[49560] = 3'b111;
        rom_memory[49561] = 3'b111;
        rom_memory[49562] = 3'b111;
        rom_memory[49563] = 3'b110;
        rom_memory[49564] = 3'b110;
        rom_memory[49565] = 3'b110;
        rom_memory[49566] = 3'b110;
        rom_memory[49567] = 3'b110;
        rom_memory[49568] = 3'b110;
        rom_memory[49569] = 3'b110;
        rom_memory[49570] = 3'b110;
        rom_memory[49571] = 3'b110;
        rom_memory[49572] = 3'b110;
        rom_memory[49573] = 3'b110;
        rom_memory[49574] = 3'b110;
        rom_memory[49575] = 3'b110;
        rom_memory[49576] = 3'b110;
        rom_memory[49577] = 3'b110;
        rom_memory[49578] = 3'b110;
        rom_memory[49579] = 3'b110;
        rom_memory[49580] = 3'b110;
        rom_memory[49581] = 3'b110;
        rom_memory[49582] = 3'b110;
        rom_memory[49583] = 3'b110;
        rom_memory[49584] = 3'b110;
        rom_memory[49585] = 3'b110;
        rom_memory[49586] = 3'b110;
        rom_memory[49587] = 3'b110;
        rom_memory[49588] = 3'b110;
        rom_memory[49589] = 3'b110;
        rom_memory[49590] = 3'b110;
        rom_memory[49591] = 3'b110;
        rom_memory[49592] = 3'b110;
        rom_memory[49593] = 3'b110;
        rom_memory[49594] = 3'b110;
        rom_memory[49595] = 3'b110;
        rom_memory[49596] = 3'b110;
        rom_memory[49597] = 3'b110;
        rom_memory[49598] = 3'b110;
        rom_memory[49599] = 3'b110;
        rom_memory[49600] = 3'b110;
        rom_memory[49601] = 3'b110;
        rom_memory[49602] = 3'b110;
        rom_memory[49603] = 3'b110;
        rom_memory[49604] = 3'b110;
        rom_memory[49605] = 3'b110;
        rom_memory[49606] = 3'b110;
        rom_memory[49607] = 3'b110;
        rom_memory[49608] = 3'b110;
        rom_memory[49609] = 3'b110;
        rom_memory[49610] = 3'b110;
        rom_memory[49611] = 3'b110;
        rom_memory[49612] = 3'b110;
        rom_memory[49613] = 3'b110;
        rom_memory[49614] = 3'b110;
        rom_memory[49615] = 3'b110;
        rom_memory[49616] = 3'b110;
        rom_memory[49617] = 3'b110;
        rom_memory[49618] = 3'b110;
        rom_memory[49619] = 3'b110;
        rom_memory[49620] = 3'b110;
        rom_memory[49621] = 3'b110;
        rom_memory[49622] = 3'b110;
        rom_memory[49623] = 3'b110;
        rom_memory[49624] = 3'b110;
        rom_memory[49625] = 3'b110;
        rom_memory[49626] = 3'b110;
        rom_memory[49627] = 3'b110;
        rom_memory[49628] = 3'b110;
        rom_memory[49629] = 3'b110;
        rom_memory[49630] = 3'b110;
        rom_memory[49631] = 3'b110;
        rom_memory[49632] = 3'b110;
        rom_memory[49633] = 3'b110;
        rom_memory[49634] = 3'b110;
        rom_memory[49635] = 3'b110;
        rom_memory[49636] = 3'b110;
        rom_memory[49637] = 3'b110;
        rom_memory[49638] = 3'b110;
        rom_memory[49639] = 3'b110;
        rom_memory[49640] = 3'b110;
        rom_memory[49641] = 3'b110;
        rom_memory[49642] = 3'b110;
        rom_memory[49643] = 3'b110;
        rom_memory[49644] = 3'b110;
        rom_memory[49645] = 3'b110;
        rom_memory[49646] = 3'b110;
        rom_memory[49647] = 3'b110;
        rom_memory[49648] = 3'b110;
        rom_memory[49649] = 3'b110;
        rom_memory[49650] = 3'b110;
        rom_memory[49651] = 3'b110;
        rom_memory[49652] = 3'b110;
        rom_memory[49653] = 3'b110;
        rom_memory[49654] = 3'b110;
        rom_memory[49655] = 3'b110;
        rom_memory[49656] = 3'b110;
        rom_memory[49657] = 3'b110;
        rom_memory[49658] = 3'b110;
        rom_memory[49659] = 3'b110;
        rom_memory[49660] = 3'b110;
        rom_memory[49661] = 3'b110;
        rom_memory[49662] = 3'b110;
        rom_memory[49663] = 3'b110;
        rom_memory[49664] = 3'b110;
        rom_memory[49665] = 3'b110;
        rom_memory[49666] = 3'b110;
        rom_memory[49667] = 3'b110;
        rom_memory[49668] = 3'b110;
        rom_memory[49669] = 3'b110;
        rom_memory[49670] = 3'b110;
        rom_memory[49671] = 3'b110;
        rom_memory[49672] = 3'b110;
        rom_memory[49673] = 3'b110;
        rom_memory[49674] = 3'b110;
        rom_memory[49675] = 3'b110;
        rom_memory[49676] = 3'b110;
        rom_memory[49677] = 3'b110;
        rom_memory[49678] = 3'b110;
        rom_memory[49679] = 3'b110;
        rom_memory[49680] = 3'b110;
        rom_memory[49681] = 3'b110;
        rom_memory[49682] = 3'b110;
        rom_memory[49683] = 3'b110;
        rom_memory[49684] = 3'b110;
        rom_memory[49685] = 3'b110;
        rom_memory[49686] = 3'b110;
        rom_memory[49687] = 3'b110;
        rom_memory[49688] = 3'b110;
        rom_memory[49689] = 3'b110;
        rom_memory[49690] = 3'b110;
        rom_memory[49691] = 3'b110;
        rom_memory[49692] = 3'b110;
        rom_memory[49693] = 3'b110;
        rom_memory[49694] = 3'b110;
        rom_memory[49695] = 3'b110;
        rom_memory[49696] = 3'b110;
        rom_memory[49697] = 3'b110;
        rom_memory[49698] = 3'b110;
        rom_memory[49699] = 3'b110;
        rom_memory[49700] = 3'b110;
        rom_memory[49701] = 3'b110;
        rom_memory[49702] = 3'b110;
        rom_memory[49703] = 3'b110;
        rom_memory[49704] = 3'b110;
        rom_memory[49705] = 3'b110;
        rom_memory[49706] = 3'b110;
        rom_memory[49707] = 3'b110;
        rom_memory[49708] = 3'b110;
        rom_memory[49709] = 3'b110;
        rom_memory[49710] = 3'b110;
        rom_memory[49711] = 3'b110;
        rom_memory[49712] = 3'b110;
        rom_memory[49713] = 3'b110;
        rom_memory[49714] = 3'b110;
        rom_memory[49715] = 3'b110;
        rom_memory[49716] = 3'b110;
        rom_memory[49717] = 3'b110;
        rom_memory[49718] = 3'b110;
        rom_memory[49719] = 3'b110;
        rom_memory[49720] = 3'b110;
        rom_memory[49721] = 3'b110;
        rom_memory[49722] = 3'b110;
        rom_memory[49723] = 3'b110;
        rom_memory[49724] = 3'b110;
        rom_memory[49725] = 3'b110;
        rom_memory[49726] = 3'b111;
        rom_memory[49727] = 3'b111;
        rom_memory[49728] = 3'b111;
        rom_memory[49729] = 3'b111;
        rom_memory[49730] = 3'b110;
        rom_memory[49731] = 3'b110;
        rom_memory[49732] = 3'b110;
        rom_memory[49733] = 3'b010;
        rom_memory[49734] = 3'b110;
        rom_memory[49735] = 3'b110;
        rom_memory[49736] = 3'b110;
        rom_memory[49737] = 3'b111;
        rom_memory[49738] = 3'b110;
        rom_memory[49739] = 3'b110;
        rom_memory[49740] = 3'b111;
        rom_memory[49741] = 3'b111;
        rom_memory[49742] = 3'b111;
        rom_memory[49743] = 3'b111;
        rom_memory[49744] = 3'b111;
        rom_memory[49745] = 3'b111;
        rom_memory[49746] = 3'b111;
        rom_memory[49747] = 3'b111;
        rom_memory[49748] = 3'b000;
        rom_memory[49749] = 3'b111;
        rom_memory[49750] = 3'b111;
        rom_memory[49751] = 3'b110;
        rom_memory[49752] = 3'b000;
        rom_memory[49753] = 3'b000;
        rom_memory[49754] = 3'b000;
        rom_memory[49755] = 3'b000;
        rom_memory[49756] = 3'b000;
        rom_memory[49757] = 3'b000;
        rom_memory[49758] = 3'b000;
        rom_memory[49759] = 3'b000;
        rom_memory[49760] = 3'b000;
        rom_memory[49761] = 3'b000;
        rom_memory[49762] = 3'b000;
        rom_memory[49763] = 3'b000;
        rom_memory[49764] = 3'b000;
        rom_memory[49765] = 3'b110;
        rom_memory[49766] = 3'b111;
        rom_memory[49767] = 3'b111;
        rom_memory[49768] = 3'b110;
        rom_memory[49769] = 3'b111;
        rom_memory[49770] = 3'b110;
        rom_memory[49771] = 3'b100;
        rom_memory[49772] = 3'b100;
        rom_memory[49773] = 3'b100;
        rom_memory[49774] = 3'b110;
        rom_memory[49775] = 3'b110;
        rom_memory[49776] = 3'b110;
        rom_memory[49777] = 3'b110;
        rom_memory[49778] = 3'b110;
        rom_memory[49779] = 3'b110;
        rom_memory[49780] = 3'b110;
        rom_memory[49781] = 3'b110;
        rom_memory[49782] = 3'b110;
        rom_memory[49783] = 3'b110;
        rom_memory[49784] = 3'b110;
        rom_memory[49785] = 3'b111;
        rom_memory[49786] = 3'b111;
        rom_memory[49787] = 3'b110;
        rom_memory[49788] = 3'b100;
        rom_memory[49789] = 3'b000;
        rom_memory[49790] = 3'b000;
        rom_memory[49791] = 3'b000;
        rom_memory[49792] = 3'b000;
        rom_memory[49793] = 3'b000;
        rom_memory[49794] = 3'b100;
        rom_memory[49795] = 3'b111;
        rom_memory[49796] = 3'b111;
        rom_memory[49797] = 3'b111;
        rom_memory[49798] = 3'b111;
        rom_memory[49799] = 3'b111;
        rom_memory[49800] = 3'b111;
        rom_memory[49801] = 3'b111;
        rom_memory[49802] = 3'b111;
        rom_memory[49803] = 3'b111;
        rom_memory[49804] = 3'b110;
        rom_memory[49805] = 3'b110;
        rom_memory[49806] = 3'b110;
        rom_memory[49807] = 3'b110;
        rom_memory[49808] = 3'b110;
        rom_memory[49809] = 3'b110;
        rom_memory[49810] = 3'b110;
        rom_memory[49811] = 3'b110;
        rom_memory[49812] = 3'b110;
        rom_memory[49813] = 3'b110;
        rom_memory[49814] = 3'b110;
        rom_memory[49815] = 3'b110;
        rom_memory[49816] = 3'b110;
        rom_memory[49817] = 3'b110;
        rom_memory[49818] = 3'b110;
        rom_memory[49819] = 3'b110;
        rom_memory[49820] = 3'b110;
        rom_memory[49821] = 3'b110;
        rom_memory[49822] = 3'b110;
        rom_memory[49823] = 3'b110;
        rom_memory[49824] = 3'b110;
        rom_memory[49825] = 3'b110;
        rom_memory[49826] = 3'b110;
        rom_memory[49827] = 3'b110;
        rom_memory[49828] = 3'b110;
        rom_memory[49829] = 3'b110;
        rom_memory[49830] = 3'b110;
        rom_memory[49831] = 3'b110;
        rom_memory[49832] = 3'b110;
        rom_memory[49833] = 3'b110;
        rom_memory[49834] = 3'b110;
        rom_memory[49835] = 3'b110;
        rom_memory[49836] = 3'b110;
        rom_memory[49837] = 3'b110;
        rom_memory[49838] = 3'b110;
        rom_memory[49839] = 3'b110;
        rom_memory[49840] = 3'b110;
        rom_memory[49841] = 3'b110;
        rom_memory[49842] = 3'b110;
        rom_memory[49843] = 3'b110;
        rom_memory[49844] = 3'b110;
        rom_memory[49845] = 3'b110;
        rom_memory[49846] = 3'b110;
        rom_memory[49847] = 3'b110;
        rom_memory[49848] = 3'b110;
        rom_memory[49849] = 3'b110;
        rom_memory[49850] = 3'b110;
        rom_memory[49851] = 3'b110;
        rom_memory[49852] = 3'b110;
        rom_memory[49853] = 3'b110;
        rom_memory[49854] = 3'b110;
        rom_memory[49855] = 3'b110;
        rom_memory[49856] = 3'b110;
        rom_memory[49857] = 3'b110;
        rom_memory[49858] = 3'b110;
        rom_memory[49859] = 3'b110;
        rom_memory[49860] = 3'b110;
        rom_memory[49861] = 3'b110;
        rom_memory[49862] = 3'b110;
        rom_memory[49863] = 3'b110;
        rom_memory[49864] = 3'b110;
        rom_memory[49865] = 3'b110;
        rom_memory[49866] = 3'b110;
        rom_memory[49867] = 3'b110;
        rom_memory[49868] = 3'b110;
        rom_memory[49869] = 3'b110;
        rom_memory[49870] = 3'b110;
        rom_memory[49871] = 3'b110;
        rom_memory[49872] = 3'b110;
        rom_memory[49873] = 3'b110;
        rom_memory[49874] = 3'b110;
        rom_memory[49875] = 3'b110;
        rom_memory[49876] = 3'b110;
        rom_memory[49877] = 3'b110;
        rom_memory[49878] = 3'b110;
        rom_memory[49879] = 3'b110;
        rom_memory[49880] = 3'b110;
        rom_memory[49881] = 3'b110;
        rom_memory[49882] = 3'b110;
        rom_memory[49883] = 3'b110;
        rom_memory[49884] = 3'b110;
        rom_memory[49885] = 3'b110;
        rom_memory[49886] = 3'b110;
        rom_memory[49887] = 3'b110;
        rom_memory[49888] = 3'b110;
        rom_memory[49889] = 3'b110;
        rom_memory[49890] = 3'b110;
        rom_memory[49891] = 3'b110;
        rom_memory[49892] = 3'b110;
        rom_memory[49893] = 3'b110;
        rom_memory[49894] = 3'b110;
        rom_memory[49895] = 3'b110;
        rom_memory[49896] = 3'b110;
        rom_memory[49897] = 3'b110;
        rom_memory[49898] = 3'b110;
        rom_memory[49899] = 3'b110;
        rom_memory[49900] = 3'b110;
        rom_memory[49901] = 3'b110;
        rom_memory[49902] = 3'b110;
        rom_memory[49903] = 3'b110;
        rom_memory[49904] = 3'b110;
        rom_memory[49905] = 3'b110;
        rom_memory[49906] = 3'b110;
        rom_memory[49907] = 3'b110;
        rom_memory[49908] = 3'b110;
        rom_memory[49909] = 3'b110;
        rom_memory[49910] = 3'b110;
        rom_memory[49911] = 3'b110;
        rom_memory[49912] = 3'b110;
        rom_memory[49913] = 3'b110;
        rom_memory[49914] = 3'b110;
        rom_memory[49915] = 3'b110;
        rom_memory[49916] = 3'b110;
        rom_memory[49917] = 3'b110;
        rom_memory[49918] = 3'b110;
        rom_memory[49919] = 3'b110;
        rom_memory[49920] = 3'b110;
        rom_memory[49921] = 3'b110;
        rom_memory[49922] = 3'b110;
        rom_memory[49923] = 3'b110;
        rom_memory[49924] = 3'b110;
        rom_memory[49925] = 3'b110;
        rom_memory[49926] = 3'b110;
        rom_memory[49927] = 3'b110;
        rom_memory[49928] = 3'b110;
        rom_memory[49929] = 3'b110;
        rom_memory[49930] = 3'b110;
        rom_memory[49931] = 3'b110;
        rom_memory[49932] = 3'b110;
        rom_memory[49933] = 3'b110;
        rom_memory[49934] = 3'b110;
        rom_memory[49935] = 3'b110;
        rom_memory[49936] = 3'b110;
        rom_memory[49937] = 3'b110;
        rom_memory[49938] = 3'b110;
        rom_memory[49939] = 3'b110;
        rom_memory[49940] = 3'b110;
        rom_memory[49941] = 3'b110;
        rom_memory[49942] = 3'b110;
        rom_memory[49943] = 3'b110;
        rom_memory[49944] = 3'b110;
        rom_memory[49945] = 3'b110;
        rom_memory[49946] = 3'b110;
        rom_memory[49947] = 3'b110;
        rom_memory[49948] = 3'b110;
        rom_memory[49949] = 3'b110;
        rom_memory[49950] = 3'b110;
        rom_memory[49951] = 3'b110;
        rom_memory[49952] = 3'b110;
        rom_memory[49953] = 3'b110;
        rom_memory[49954] = 3'b110;
        rom_memory[49955] = 3'b110;
        rom_memory[49956] = 3'b110;
        rom_memory[49957] = 3'b110;
        rom_memory[49958] = 3'b110;
        rom_memory[49959] = 3'b110;
        rom_memory[49960] = 3'b110;
        rom_memory[49961] = 3'b110;
        rom_memory[49962] = 3'b110;
        rom_memory[49963] = 3'b110;
        rom_memory[49964] = 3'b110;
        rom_memory[49965] = 3'b110;
        rom_memory[49966] = 3'b111;
        rom_memory[49967] = 3'b111;
        rom_memory[49968] = 3'b111;
        rom_memory[49969] = 3'b111;
        rom_memory[49970] = 3'b010;
        rom_memory[49971] = 3'b000;
        rom_memory[49972] = 3'b110;
        rom_memory[49973] = 3'b110;
        rom_memory[49974] = 3'b110;
        rom_memory[49975] = 3'b110;
        rom_memory[49976] = 3'b111;
        rom_memory[49977] = 3'b111;
        rom_memory[49978] = 3'b110;
        rom_memory[49979] = 3'b111;
        rom_memory[49980] = 3'b111;
        rom_memory[49981] = 3'b111;
        rom_memory[49982] = 3'b111;
        rom_memory[49983] = 3'b111;
        rom_memory[49984] = 3'b111;
        rom_memory[49985] = 3'b111;
        rom_memory[49986] = 3'b111;
        rom_memory[49987] = 3'b111;
        rom_memory[49988] = 3'b111;
        rom_memory[49989] = 3'b111;
        rom_memory[49990] = 3'b111;
        rom_memory[49991] = 3'b111;
        rom_memory[49992] = 3'b111;
        rom_memory[49993] = 3'b000;
        rom_memory[49994] = 3'b000;
        rom_memory[49995] = 3'b000;
        rom_memory[49996] = 3'b000;
        rom_memory[49997] = 3'b000;
        rom_memory[49998] = 3'b000;
        rom_memory[49999] = 3'b000;
        rom_memory[50000] = 3'b000;
        rom_memory[50001] = 3'b000;
        rom_memory[50002] = 3'b000;
        rom_memory[50003] = 3'b000;
        rom_memory[50004] = 3'b000;
        rom_memory[50005] = 3'b111;
        rom_memory[50006] = 3'b111;
        rom_memory[50007] = 3'b111;
        rom_memory[50008] = 3'b110;
        rom_memory[50009] = 3'b111;
        rom_memory[50010] = 3'b110;
        rom_memory[50011] = 3'b100;
        rom_memory[50012] = 3'b100;
        rom_memory[50013] = 3'b100;
        rom_memory[50014] = 3'b110;
        rom_memory[50015] = 3'b110;
        rom_memory[50016] = 3'b110;
        rom_memory[50017] = 3'b110;
        rom_memory[50018] = 3'b110;
        rom_memory[50019] = 3'b110;
        rom_memory[50020] = 3'b110;
        rom_memory[50021] = 3'b110;
        rom_memory[50022] = 3'b110;
        rom_memory[50023] = 3'b110;
        rom_memory[50024] = 3'b111;
        rom_memory[50025] = 3'b111;
        rom_memory[50026] = 3'b111;
        rom_memory[50027] = 3'b111;
        rom_memory[50028] = 3'b100;
        rom_memory[50029] = 3'b000;
        rom_memory[50030] = 3'b000;
        rom_memory[50031] = 3'b000;
        rom_memory[50032] = 3'b000;
        rom_memory[50033] = 3'b000;
        rom_memory[50034] = 3'b100;
        rom_memory[50035] = 3'b111;
        rom_memory[50036] = 3'b111;
        rom_memory[50037] = 3'b111;
        rom_memory[50038] = 3'b111;
        rom_memory[50039] = 3'b111;
        rom_memory[50040] = 3'b111;
        rom_memory[50041] = 3'b111;
        rom_memory[50042] = 3'b111;
        rom_memory[50043] = 3'b111;
        rom_memory[50044] = 3'b110;
        rom_memory[50045] = 3'b110;
        rom_memory[50046] = 3'b110;
        rom_memory[50047] = 3'b110;
        rom_memory[50048] = 3'b110;
        rom_memory[50049] = 3'b110;
        rom_memory[50050] = 3'b110;
        rom_memory[50051] = 3'b110;
        rom_memory[50052] = 3'b110;
        rom_memory[50053] = 3'b110;
        rom_memory[50054] = 3'b110;
        rom_memory[50055] = 3'b110;
        rom_memory[50056] = 3'b110;
        rom_memory[50057] = 3'b110;
        rom_memory[50058] = 3'b110;
        rom_memory[50059] = 3'b110;
        rom_memory[50060] = 3'b110;
        rom_memory[50061] = 3'b110;
        rom_memory[50062] = 3'b110;
        rom_memory[50063] = 3'b110;
        rom_memory[50064] = 3'b110;
        rom_memory[50065] = 3'b110;
        rom_memory[50066] = 3'b110;
        rom_memory[50067] = 3'b110;
        rom_memory[50068] = 3'b110;
        rom_memory[50069] = 3'b110;
        rom_memory[50070] = 3'b110;
        rom_memory[50071] = 3'b110;
        rom_memory[50072] = 3'b110;
        rom_memory[50073] = 3'b110;
        rom_memory[50074] = 3'b110;
        rom_memory[50075] = 3'b110;
        rom_memory[50076] = 3'b110;
        rom_memory[50077] = 3'b110;
        rom_memory[50078] = 3'b110;
        rom_memory[50079] = 3'b110;
        rom_memory[50080] = 3'b110;
        rom_memory[50081] = 3'b110;
        rom_memory[50082] = 3'b110;
        rom_memory[50083] = 3'b110;
        rom_memory[50084] = 3'b110;
        rom_memory[50085] = 3'b110;
        rom_memory[50086] = 3'b110;
        rom_memory[50087] = 3'b110;
        rom_memory[50088] = 3'b110;
        rom_memory[50089] = 3'b110;
        rom_memory[50090] = 3'b110;
        rom_memory[50091] = 3'b110;
        rom_memory[50092] = 3'b110;
        rom_memory[50093] = 3'b110;
        rom_memory[50094] = 3'b110;
        rom_memory[50095] = 3'b110;
        rom_memory[50096] = 3'b110;
        rom_memory[50097] = 3'b110;
        rom_memory[50098] = 3'b110;
        rom_memory[50099] = 3'b110;
        rom_memory[50100] = 3'b110;
        rom_memory[50101] = 3'b110;
        rom_memory[50102] = 3'b110;
        rom_memory[50103] = 3'b110;
        rom_memory[50104] = 3'b110;
        rom_memory[50105] = 3'b110;
        rom_memory[50106] = 3'b110;
        rom_memory[50107] = 3'b110;
        rom_memory[50108] = 3'b110;
        rom_memory[50109] = 3'b110;
        rom_memory[50110] = 3'b110;
        rom_memory[50111] = 3'b110;
        rom_memory[50112] = 3'b110;
        rom_memory[50113] = 3'b110;
        rom_memory[50114] = 3'b110;
        rom_memory[50115] = 3'b110;
        rom_memory[50116] = 3'b110;
        rom_memory[50117] = 3'b110;
        rom_memory[50118] = 3'b110;
        rom_memory[50119] = 3'b110;
        rom_memory[50120] = 3'b110;
        rom_memory[50121] = 3'b110;
        rom_memory[50122] = 3'b110;
        rom_memory[50123] = 3'b110;
        rom_memory[50124] = 3'b110;
        rom_memory[50125] = 3'b110;
        rom_memory[50126] = 3'b110;
        rom_memory[50127] = 3'b110;
        rom_memory[50128] = 3'b110;
        rom_memory[50129] = 3'b110;
        rom_memory[50130] = 3'b110;
        rom_memory[50131] = 3'b110;
        rom_memory[50132] = 3'b110;
        rom_memory[50133] = 3'b110;
        rom_memory[50134] = 3'b110;
        rom_memory[50135] = 3'b110;
        rom_memory[50136] = 3'b110;
        rom_memory[50137] = 3'b110;
        rom_memory[50138] = 3'b110;
        rom_memory[50139] = 3'b110;
        rom_memory[50140] = 3'b110;
        rom_memory[50141] = 3'b110;
        rom_memory[50142] = 3'b110;
        rom_memory[50143] = 3'b110;
        rom_memory[50144] = 3'b110;
        rom_memory[50145] = 3'b110;
        rom_memory[50146] = 3'b110;
        rom_memory[50147] = 3'b110;
        rom_memory[50148] = 3'b110;
        rom_memory[50149] = 3'b110;
        rom_memory[50150] = 3'b110;
        rom_memory[50151] = 3'b110;
        rom_memory[50152] = 3'b110;
        rom_memory[50153] = 3'b110;
        rom_memory[50154] = 3'b110;
        rom_memory[50155] = 3'b110;
        rom_memory[50156] = 3'b110;
        rom_memory[50157] = 3'b110;
        rom_memory[50158] = 3'b110;
        rom_memory[50159] = 3'b110;
        rom_memory[50160] = 3'b111;
        rom_memory[50161] = 3'b111;
        rom_memory[50162] = 3'b110;
        rom_memory[50163] = 3'b110;
        rom_memory[50164] = 3'b110;
        rom_memory[50165] = 3'b110;
        rom_memory[50166] = 3'b110;
        rom_memory[50167] = 3'b110;
        rom_memory[50168] = 3'b110;
        rom_memory[50169] = 3'b110;
        rom_memory[50170] = 3'b110;
        rom_memory[50171] = 3'b110;
        rom_memory[50172] = 3'b110;
        rom_memory[50173] = 3'b110;
        rom_memory[50174] = 3'b110;
        rom_memory[50175] = 3'b110;
        rom_memory[50176] = 3'b110;
        rom_memory[50177] = 3'b110;
        rom_memory[50178] = 3'b110;
        rom_memory[50179] = 3'b100;
        rom_memory[50180] = 3'b100;
        rom_memory[50181] = 3'b100;
        rom_memory[50182] = 3'b110;
        rom_memory[50183] = 3'b110;
        rom_memory[50184] = 3'b110;
        rom_memory[50185] = 3'b110;
        rom_memory[50186] = 3'b110;
        rom_memory[50187] = 3'b110;
        rom_memory[50188] = 3'b110;
        rom_memory[50189] = 3'b110;
        rom_memory[50190] = 3'b110;
        rom_memory[50191] = 3'b110;
        rom_memory[50192] = 3'b110;
        rom_memory[50193] = 3'b110;
        rom_memory[50194] = 3'b110;
        rom_memory[50195] = 3'b110;
        rom_memory[50196] = 3'b110;
        rom_memory[50197] = 3'b110;
        rom_memory[50198] = 3'b110;
        rom_memory[50199] = 3'b110;
        rom_memory[50200] = 3'b110;
        rom_memory[50201] = 3'b110;
        rom_memory[50202] = 3'b110;
        rom_memory[50203] = 3'b110;
        rom_memory[50204] = 3'b111;
        rom_memory[50205] = 3'b111;
        rom_memory[50206] = 3'b111;
        rom_memory[50207] = 3'b111;
        rom_memory[50208] = 3'b111;
        rom_memory[50209] = 3'b111;
        rom_memory[50210] = 3'b000;
        rom_memory[50211] = 3'b000;
        rom_memory[50212] = 3'b110;
        rom_memory[50213] = 3'b110;
        rom_memory[50214] = 3'b110;
        rom_memory[50215] = 3'b111;
        rom_memory[50216] = 3'b111;
        rom_memory[50217] = 3'b111;
        rom_memory[50218] = 3'b111;
        rom_memory[50219] = 3'b111;
        rom_memory[50220] = 3'b111;
        rom_memory[50221] = 3'b111;
        rom_memory[50222] = 3'b111;
        rom_memory[50223] = 3'b111;
        rom_memory[50224] = 3'b111;
        rom_memory[50225] = 3'b111;
        rom_memory[50226] = 3'b000;
        rom_memory[50227] = 3'b100;
        rom_memory[50228] = 3'b111;
        rom_memory[50229] = 3'b111;
        rom_memory[50230] = 3'b111;
        rom_memory[50231] = 3'b111;
        rom_memory[50232] = 3'b111;
        rom_memory[50233] = 3'b000;
        rom_memory[50234] = 3'b000;
        rom_memory[50235] = 3'b000;
        rom_memory[50236] = 3'b000;
        rom_memory[50237] = 3'b000;
        rom_memory[50238] = 3'b000;
        rom_memory[50239] = 3'b000;
        rom_memory[50240] = 3'b000;
        rom_memory[50241] = 3'b000;
        rom_memory[50242] = 3'b000;
        rom_memory[50243] = 3'b000;
        rom_memory[50244] = 3'b000;
        rom_memory[50245] = 3'b111;
        rom_memory[50246] = 3'b111;
        rom_memory[50247] = 3'b111;
        rom_memory[50248] = 3'b110;
        rom_memory[50249] = 3'b111;
        rom_memory[50250] = 3'b111;
        rom_memory[50251] = 3'b000;
        rom_memory[50252] = 3'b100;
        rom_memory[50253] = 3'b110;
        rom_memory[50254] = 3'b111;
        rom_memory[50255] = 3'b100;
        rom_memory[50256] = 3'b110;
        rom_memory[50257] = 3'b110;
        rom_memory[50258] = 3'b110;
        rom_memory[50259] = 3'b110;
        rom_memory[50260] = 3'b111;
        rom_memory[50261] = 3'b111;
        rom_memory[50262] = 3'b111;
        rom_memory[50263] = 3'b111;
        rom_memory[50264] = 3'b111;
        rom_memory[50265] = 3'b111;
        rom_memory[50266] = 3'b111;
        rom_memory[50267] = 3'b111;
        rom_memory[50268] = 3'b100;
        rom_memory[50269] = 3'b000;
        rom_memory[50270] = 3'b000;
        rom_memory[50271] = 3'b000;
        rom_memory[50272] = 3'b000;
        rom_memory[50273] = 3'b000;
        rom_memory[50274] = 3'b000;
        rom_memory[50275] = 3'b100;
        rom_memory[50276] = 3'b111;
        rom_memory[50277] = 3'b111;
        rom_memory[50278] = 3'b111;
        rom_memory[50279] = 3'b111;
        rom_memory[50280] = 3'b111;
        rom_memory[50281] = 3'b111;
        rom_memory[50282] = 3'b111;
        rom_memory[50283] = 3'b111;
        rom_memory[50284] = 3'b111;
        rom_memory[50285] = 3'b110;
        rom_memory[50286] = 3'b110;
        rom_memory[50287] = 3'b110;
        rom_memory[50288] = 3'b110;
        rom_memory[50289] = 3'b110;
        rom_memory[50290] = 3'b110;
        rom_memory[50291] = 3'b110;
        rom_memory[50292] = 3'b110;
        rom_memory[50293] = 3'b110;
        rom_memory[50294] = 3'b110;
        rom_memory[50295] = 3'b110;
        rom_memory[50296] = 3'b110;
        rom_memory[50297] = 3'b110;
        rom_memory[50298] = 3'b110;
        rom_memory[50299] = 3'b110;
        rom_memory[50300] = 3'b110;
        rom_memory[50301] = 3'b110;
        rom_memory[50302] = 3'b110;
        rom_memory[50303] = 3'b110;
        rom_memory[50304] = 3'b110;
        rom_memory[50305] = 3'b110;
        rom_memory[50306] = 3'b110;
        rom_memory[50307] = 3'b110;
        rom_memory[50308] = 3'b110;
        rom_memory[50309] = 3'b110;
        rom_memory[50310] = 3'b110;
        rom_memory[50311] = 3'b110;
        rom_memory[50312] = 3'b110;
        rom_memory[50313] = 3'b110;
        rom_memory[50314] = 3'b110;
        rom_memory[50315] = 3'b110;
        rom_memory[50316] = 3'b110;
        rom_memory[50317] = 3'b110;
        rom_memory[50318] = 3'b110;
        rom_memory[50319] = 3'b110;
        rom_memory[50320] = 3'b110;
        rom_memory[50321] = 3'b110;
        rom_memory[50322] = 3'b110;
        rom_memory[50323] = 3'b110;
        rom_memory[50324] = 3'b110;
        rom_memory[50325] = 3'b110;
        rom_memory[50326] = 3'b110;
        rom_memory[50327] = 3'b110;
        rom_memory[50328] = 3'b110;
        rom_memory[50329] = 3'b110;
        rom_memory[50330] = 3'b110;
        rom_memory[50331] = 3'b110;
        rom_memory[50332] = 3'b110;
        rom_memory[50333] = 3'b110;
        rom_memory[50334] = 3'b110;
        rom_memory[50335] = 3'b110;
        rom_memory[50336] = 3'b110;
        rom_memory[50337] = 3'b110;
        rom_memory[50338] = 3'b110;
        rom_memory[50339] = 3'b110;
        rom_memory[50340] = 3'b110;
        rom_memory[50341] = 3'b110;
        rom_memory[50342] = 3'b110;
        rom_memory[50343] = 3'b110;
        rom_memory[50344] = 3'b110;
        rom_memory[50345] = 3'b110;
        rom_memory[50346] = 3'b110;
        rom_memory[50347] = 3'b110;
        rom_memory[50348] = 3'b110;
        rom_memory[50349] = 3'b110;
        rom_memory[50350] = 3'b110;
        rom_memory[50351] = 3'b110;
        rom_memory[50352] = 3'b110;
        rom_memory[50353] = 3'b110;
        rom_memory[50354] = 3'b110;
        rom_memory[50355] = 3'b110;
        rom_memory[50356] = 3'b110;
        rom_memory[50357] = 3'b110;
        rom_memory[50358] = 3'b110;
        rom_memory[50359] = 3'b110;
        rom_memory[50360] = 3'b110;
        rom_memory[50361] = 3'b110;
        rom_memory[50362] = 3'b110;
        rom_memory[50363] = 3'b110;
        rom_memory[50364] = 3'b110;
        rom_memory[50365] = 3'b110;
        rom_memory[50366] = 3'b110;
        rom_memory[50367] = 3'b110;
        rom_memory[50368] = 3'b110;
        rom_memory[50369] = 3'b110;
        rom_memory[50370] = 3'b110;
        rom_memory[50371] = 3'b110;
        rom_memory[50372] = 3'b110;
        rom_memory[50373] = 3'b110;
        rom_memory[50374] = 3'b110;
        rom_memory[50375] = 3'b110;
        rom_memory[50376] = 3'b110;
        rom_memory[50377] = 3'b110;
        rom_memory[50378] = 3'b110;
        rom_memory[50379] = 3'b110;
        rom_memory[50380] = 3'b110;
        rom_memory[50381] = 3'b110;
        rom_memory[50382] = 3'b110;
        rom_memory[50383] = 3'b110;
        rom_memory[50384] = 3'b110;
        rom_memory[50385] = 3'b110;
        rom_memory[50386] = 3'b110;
        rom_memory[50387] = 3'b110;
        rom_memory[50388] = 3'b110;
        rom_memory[50389] = 3'b110;
        rom_memory[50390] = 3'b110;
        rom_memory[50391] = 3'b110;
        rom_memory[50392] = 3'b110;
        rom_memory[50393] = 3'b110;
        rom_memory[50394] = 3'b110;
        rom_memory[50395] = 3'b110;
        rom_memory[50396] = 3'b110;
        rom_memory[50397] = 3'b110;
        rom_memory[50398] = 3'b110;
        rom_memory[50399] = 3'b110;
        rom_memory[50400] = 3'b110;
        rom_memory[50401] = 3'b110;
        rom_memory[50402] = 3'b110;
        rom_memory[50403] = 3'b110;
        rom_memory[50404] = 3'b110;
        rom_memory[50405] = 3'b110;
        rom_memory[50406] = 3'b110;
        rom_memory[50407] = 3'b110;
        rom_memory[50408] = 3'b110;
        rom_memory[50409] = 3'b110;
        rom_memory[50410] = 3'b111;
        rom_memory[50411] = 3'b110;
        rom_memory[50412] = 3'b110;
        rom_memory[50413] = 3'b110;
        rom_memory[50414] = 3'b110;
        rom_memory[50415] = 3'b110;
        rom_memory[50416] = 3'b110;
        rom_memory[50417] = 3'b110;
        rom_memory[50418] = 3'b100;
        rom_memory[50419] = 3'b100;
        rom_memory[50420] = 3'b100;
        rom_memory[50421] = 3'b100;
        rom_memory[50422] = 3'b100;
        rom_memory[50423] = 3'b100;
        rom_memory[50424] = 3'b100;
        rom_memory[50425] = 3'b100;
        rom_memory[50426] = 3'b110;
        rom_memory[50427] = 3'b110;
        rom_memory[50428] = 3'b110;
        rom_memory[50429] = 3'b110;
        rom_memory[50430] = 3'b110;
        rom_memory[50431] = 3'b110;
        rom_memory[50432] = 3'b110;
        rom_memory[50433] = 3'b110;
        rom_memory[50434] = 3'b110;
        rom_memory[50435] = 3'b110;
        rom_memory[50436] = 3'b110;
        rom_memory[50437] = 3'b110;
        rom_memory[50438] = 3'b110;
        rom_memory[50439] = 3'b110;
        rom_memory[50440] = 3'b110;
        rom_memory[50441] = 3'b110;
        rom_memory[50442] = 3'b110;
        rom_memory[50443] = 3'b110;
        rom_memory[50444] = 3'b111;
        rom_memory[50445] = 3'b111;
        rom_memory[50446] = 3'b111;
        rom_memory[50447] = 3'b111;
        rom_memory[50448] = 3'b110;
        rom_memory[50449] = 3'b110;
        rom_memory[50450] = 3'b000;
        rom_memory[50451] = 3'b000;
        rom_memory[50452] = 3'b110;
        rom_memory[50453] = 3'b110;
        rom_memory[50454] = 3'b110;
        rom_memory[50455] = 3'b110;
        rom_memory[50456] = 3'b111;
        rom_memory[50457] = 3'b111;
        rom_memory[50458] = 3'b111;
        rom_memory[50459] = 3'b111;
        rom_memory[50460] = 3'b111;
        rom_memory[50461] = 3'b111;
        rom_memory[50462] = 3'b111;
        rom_memory[50463] = 3'b111;
        rom_memory[50464] = 3'b111;
        rom_memory[50465] = 3'b111;
        rom_memory[50466] = 3'b110;
        rom_memory[50467] = 3'b100;
        rom_memory[50468] = 3'b111;
        rom_memory[50469] = 3'b111;
        rom_memory[50470] = 3'b111;
        rom_memory[50471] = 3'b111;
        rom_memory[50472] = 3'b111;
        rom_memory[50473] = 3'b111;
        rom_memory[50474] = 3'b100;
        rom_memory[50475] = 3'b000;
        rom_memory[50476] = 3'b000;
        rom_memory[50477] = 3'b000;
        rom_memory[50478] = 3'b000;
        rom_memory[50479] = 3'b000;
        rom_memory[50480] = 3'b000;
        rom_memory[50481] = 3'b000;
        rom_memory[50482] = 3'b000;
        rom_memory[50483] = 3'b000;
        rom_memory[50484] = 3'b000;
        rom_memory[50485] = 3'b111;
        rom_memory[50486] = 3'b111;
        rom_memory[50487] = 3'b111;
        rom_memory[50488] = 3'b110;
        rom_memory[50489] = 3'b111;
        rom_memory[50490] = 3'b111;
        rom_memory[50491] = 3'b111;
        rom_memory[50492] = 3'b111;
        rom_memory[50493] = 3'b111;
        rom_memory[50494] = 3'b110;
        rom_memory[50495] = 3'b100;
        rom_memory[50496] = 3'b100;
        rom_memory[50497] = 3'b110;
        rom_memory[50498] = 3'b110;
        rom_memory[50499] = 3'b110;
        rom_memory[50500] = 3'b111;
        rom_memory[50501] = 3'b111;
        rom_memory[50502] = 3'b111;
        rom_memory[50503] = 3'b111;
        rom_memory[50504] = 3'b111;
        rom_memory[50505] = 3'b111;
        rom_memory[50506] = 3'b111;
        rom_memory[50507] = 3'b111;
        rom_memory[50508] = 3'b100;
        rom_memory[50509] = 3'b000;
        rom_memory[50510] = 3'b000;
        rom_memory[50511] = 3'b000;
        rom_memory[50512] = 3'b000;
        rom_memory[50513] = 3'b000;
        rom_memory[50514] = 3'b000;
        rom_memory[50515] = 3'b000;
        rom_memory[50516] = 3'b100;
        rom_memory[50517] = 3'b111;
        rom_memory[50518] = 3'b111;
        rom_memory[50519] = 3'b111;
        rom_memory[50520] = 3'b111;
        rom_memory[50521] = 3'b111;
        rom_memory[50522] = 3'b111;
        rom_memory[50523] = 3'b111;
        rom_memory[50524] = 3'b111;
        rom_memory[50525] = 3'b110;
        rom_memory[50526] = 3'b110;
        rom_memory[50527] = 3'b110;
        rom_memory[50528] = 3'b110;
        rom_memory[50529] = 3'b110;
        rom_memory[50530] = 3'b110;
        rom_memory[50531] = 3'b110;
        rom_memory[50532] = 3'b110;
        rom_memory[50533] = 3'b110;
        rom_memory[50534] = 3'b110;
        rom_memory[50535] = 3'b110;
        rom_memory[50536] = 3'b110;
        rom_memory[50537] = 3'b110;
        rom_memory[50538] = 3'b110;
        rom_memory[50539] = 3'b110;
        rom_memory[50540] = 3'b110;
        rom_memory[50541] = 3'b110;
        rom_memory[50542] = 3'b110;
        rom_memory[50543] = 3'b110;
        rom_memory[50544] = 3'b110;
        rom_memory[50545] = 3'b110;
        rom_memory[50546] = 3'b110;
        rom_memory[50547] = 3'b110;
        rom_memory[50548] = 3'b110;
        rom_memory[50549] = 3'b110;
        rom_memory[50550] = 3'b110;
        rom_memory[50551] = 3'b110;
        rom_memory[50552] = 3'b110;
        rom_memory[50553] = 3'b110;
        rom_memory[50554] = 3'b110;
        rom_memory[50555] = 3'b110;
        rom_memory[50556] = 3'b110;
        rom_memory[50557] = 3'b110;
        rom_memory[50558] = 3'b110;
        rom_memory[50559] = 3'b110;
        rom_memory[50560] = 3'b110;
        rom_memory[50561] = 3'b110;
        rom_memory[50562] = 3'b110;
        rom_memory[50563] = 3'b110;
        rom_memory[50564] = 3'b110;
        rom_memory[50565] = 3'b110;
        rom_memory[50566] = 3'b110;
        rom_memory[50567] = 3'b110;
        rom_memory[50568] = 3'b110;
        rom_memory[50569] = 3'b110;
        rom_memory[50570] = 3'b110;
        rom_memory[50571] = 3'b110;
        rom_memory[50572] = 3'b110;
        rom_memory[50573] = 3'b110;
        rom_memory[50574] = 3'b110;
        rom_memory[50575] = 3'b110;
        rom_memory[50576] = 3'b110;
        rom_memory[50577] = 3'b110;
        rom_memory[50578] = 3'b110;
        rom_memory[50579] = 3'b110;
        rom_memory[50580] = 3'b110;
        rom_memory[50581] = 3'b110;
        rom_memory[50582] = 3'b110;
        rom_memory[50583] = 3'b110;
        rom_memory[50584] = 3'b110;
        rom_memory[50585] = 3'b110;
        rom_memory[50586] = 3'b110;
        rom_memory[50587] = 3'b110;
        rom_memory[50588] = 3'b110;
        rom_memory[50589] = 3'b110;
        rom_memory[50590] = 3'b110;
        rom_memory[50591] = 3'b110;
        rom_memory[50592] = 3'b110;
        rom_memory[50593] = 3'b110;
        rom_memory[50594] = 3'b110;
        rom_memory[50595] = 3'b110;
        rom_memory[50596] = 3'b110;
        rom_memory[50597] = 3'b110;
        rom_memory[50598] = 3'b110;
        rom_memory[50599] = 3'b110;
        rom_memory[50600] = 3'b110;
        rom_memory[50601] = 3'b110;
        rom_memory[50602] = 3'b110;
        rom_memory[50603] = 3'b110;
        rom_memory[50604] = 3'b110;
        rom_memory[50605] = 3'b110;
        rom_memory[50606] = 3'b110;
        rom_memory[50607] = 3'b110;
        rom_memory[50608] = 3'b110;
        rom_memory[50609] = 3'b110;
        rom_memory[50610] = 3'b110;
        rom_memory[50611] = 3'b110;
        rom_memory[50612] = 3'b110;
        rom_memory[50613] = 3'b110;
        rom_memory[50614] = 3'b110;
        rom_memory[50615] = 3'b110;
        rom_memory[50616] = 3'b110;
        rom_memory[50617] = 3'b110;
        rom_memory[50618] = 3'b110;
        rom_memory[50619] = 3'b110;
        rom_memory[50620] = 3'b110;
        rom_memory[50621] = 3'b110;
        rom_memory[50622] = 3'b110;
        rom_memory[50623] = 3'b110;
        rom_memory[50624] = 3'b110;
        rom_memory[50625] = 3'b110;
        rom_memory[50626] = 3'b110;
        rom_memory[50627] = 3'b110;
        rom_memory[50628] = 3'b110;
        rom_memory[50629] = 3'b110;
        rom_memory[50630] = 3'b110;
        rom_memory[50631] = 3'b110;
        rom_memory[50632] = 3'b110;
        rom_memory[50633] = 3'b110;
        rom_memory[50634] = 3'b110;
        rom_memory[50635] = 3'b110;
        rom_memory[50636] = 3'b110;
        rom_memory[50637] = 3'b110;
        rom_memory[50638] = 3'b110;
        rom_memory[50639] = 3'b110;
        rom_memory[50640] = 3'b110;
        rom_memory[50641] = 3'b110;
        rom_memory[50642] = 3'b110;
        rom_memory[50643] = 3'b110;
        rom_memory[50644] = 3'b110;
        rom_memory[50645] = 3'b110;
        rom_memory[50646] = 3'b110;
        rom_memory[50647] = 3'b110;
        rom_memory[50648] = 3'b110;
        rom_memory[50649] = 3'b110;
        rom_memory[50650] = 3'b111;
        rom_memory[50651] = 3'b111;
        rom_memory[50652] = 3'b110;
        rom_memory[50653] = 3'b110;
        rom_memory[50654] = 3'b110;
        rom_memory[50655] = 3'b110;
        rom_memory[50656] = 3'b110;
        rom_memory[50657] = 3'b110;
        rom_memory[50658] = 3'b100;
        rom_memory[50659] = 3'b100;
        rom_memory[50660] = 3'b100;
        rom_memory[50661] = 3'b100;
        rom_memory[50662] = 3'b100;
        rom_memory[50663] = 3'b100;
        rom_memory[50664] = 3'b100;
        rom_memory[50665] = 3'b100;
        rom_memory[50666] = 3'b110;
        rom_memory[50667] = 3'b110;
        rom_memory[50668] = 3'b110;
        rom_memory[50669] = 3'b110;
        rom_memory[50670] = 3'b110;
        rom_memory[50671] = 3'b110;
        rom_memory[50672] = 3'b110;
        rom_memory[50673] = 3'b110;
        rom_memory[50674] = 3'b110;
        rom_memory[50675] = 3'b110;
        rom_memory[50676] = 3'b110;
        rom_memory[50677] = 3'b110;
        rom_memory[50678] = 3'b110;
        rom_memory[50679] = 3'b110;
        rom_memory[50680] = 3'b110;
        rom_memory[50681] = 3'b110;
        rom_memory[50682] = 3'b110;
        rom_memory[50683] = 3'b110;
        rom_memory[50684] = 3'b111;
        rom_memory[50685] = 3'b111;
        rom_memory[50686] = 3'b111;
        rom_memory[50687] = 3'b111;
        rom_memory[50688] = 3'b110;
        rom_memory[50689] = 3'b100;
        rom_memory[50690] = 3'b100;
        rom_memory[50691] = 3'b000;
        rom_memory[50692] = 3'b000;
        rom_memory[50693] = 3'b100;
        rom_memory[50694] = 3'b110;
        rom_memory[50695] = 3'b111;
        rom_memory[50696] = 3'b111;
        rom_memory[50697] = 3'b111;
        rom_memory[50698] = 3'b111;
        rom_memory[50699] = 3'b111;
        rom_memory[50700] = 3'b111;
        rom_memory[50701] = 3'b111;
        rom_memory[50702] = 3'b111;
        rom_memory[50703] = 3'b111;
        rom_memory[50704] = 3'b111;
        rom_memory[50705] = 3'b111;
        rom_memory[50706] = 3'b100;
        rom_memory[50707] = 3'b111;
        rom_memory[50708] = 3'b111;
        rom_memory[50709] = 3'b111;
        rom_memory[50710] = 3'b111;
        rom_memory[50711] = 3'b111;
        rom_memory[50712] = 3'b111;
        rom_memory[50713] = 3'b110;
        rom_memory[50714] = 3'b000;
        rom_memory[50715] = 3'b000;
        rom_memory[50716] = 3'b000;
        rom_memory[50717] = 3'b000;
        rom_memory[50718] = 3'b000;
        rom_memory[50719] = 3'b000;
        rom_memory[50720] = 3'b000;
        rom_memory[50721] = 3'b000;
        rom_memory[50722] = 3'b000;
        rom_memory[50723] = 3'b000;
        rom_memory[50724] = 3'b000;
        rom_memory[50725] = 3'b111;
        rom_memory[50726] = 3'b111;
        rom_memory[50727] = 3'b111;
        rom_memory[50728] = 3'b110;
        rom_memory[50729] = 3'b111;
        rom_memory[50730] = 3'b111;
        rom_memory[50731] = 3'b111;
        rom_memory[50732] = 3'b111;
        rom_memory[50733] = 3'b111;
        rom_memory[50734] = 3'b110;
        rom_memory[50735] = 3'b000;
        rom_memory[50736] = 3'b100;
        rom_memory[50737] = 3'b100;
        rom_memory[50738] = 3'b110;
        rom_memory[50739] = 3'b110;
        rom_memory[50740] = 3'b111;
        rom_memory[50741] = 3'b111;
        rom_memory[50742] = 3'b111;
        rom_memory[50743] = 3'b111;
        rom_memory[50744] = 3'b111;
        rom_memory[50745] = 3'b111;
        rom_memory[50746] = 3'b111;
        rom_memory[50747] = 3'b111;
        rom_memory[50748] = 3'b100;
        rom_memory[50749] = 3'b100;
        rom_memory[50750] = 3'b000;
        rom_memory[50751] = 3'b000;
        rom_memory[50752] = 3'b000;
        rom_memory[50753] = 3'b000;
        rom_memory[50754] = 3'b000;
        rom_memory[50755] = 3'b000;
        rom_memory[50756] = 3'b100;
        rom_memory[50757] = 3'b101;
        rom_memory[50758] = 3'b111;
        rom_memory[50759] = 3'b111;
        rom_memory[50760] = 3'b111;
        rom_memory[50761] = 3'b111;
        rom_memory[50762] = 3'b111;
        rom_memory[50763] = 3'b111;
        rom_memory[50764] = 3'b111;
        rom_memory[50765] = 3'b110;
        rom_memory[50766] = 3'b110;
        rom_memory[50767] = 3'b110;
        rom_memory[50768] = 3'b110;
        rom_memory[50769] = 3'b110;
        rom_memory[50770] = 3'b110;
        rom_memory[50771] = 3'b110;
        rom_memory[50772] = 3'b110;
        rom_memory[50773] = 3'b110;
        rom_memory[50774] = 3'b110;
        rom_memory[50775] = 3'b110;
        rom_memory[50776] = 3'b110;
        rom_memory[50777] = 3'b110;
        rom_memory[50778] = 3'b110;
        rom_memory[50779] = 3'b110;
        rom_memory[50780] = 3'b110;
        rom_memory[50781] = 3'b110;
        rom_memory[50782] = 3'b110;
        rom_memory[50783] = 3'b110;
        rom_memory[50784] = 3'b110;
        rom_memory[50785] = 3'b110;
        rom_memory[50786] = 3'b110;
        rom_memory[50787] = 3'b110;
        rom_memory[50788] = 3'b110;
        rom_memory[50789] = 3'b110;
        rom_memory[50790] = 3'b110;
        rom_memory[50791] = 3'b110;
        rom_memory[50792] = 3'b110;
        rom_memory[50793] = 3'b110;
        rom_memory[50794] = 3'b110;
        rom_memory[50795] = 3'b110;
        rom_memory[50796] = 3'b110;
        rom_memory[50797] = 3'b110;
        rom_memory[50798] = 3'b110;
        rom_memory[50799] = 3'b110;
        rom_memory[50800] = 3'b110;
        rom_memory[50801] = 3'b110;
        rom_memory[50802] = 3'b110;
        rom_memory[50803] = 3'b110;
        rom_memory[50804] = 3'b110;
        rom_memory[50805] = 3'b110;
        rom_memory[50806] = 3'b110;
        rom_memory[50807] = 3'b110;
        rom_memory[50808] = 3'b110;
        rom_memory[50809] = 3'b110;
        rom_memory[50810] = 3'b110;
        rom_memory[50811] = 3'b110;
        rom_memory[50812] = 3'b110;
        rom_memory[50813] = 3'b110;
        rom_memory[50814] = 3'b110;
        rom_memory[50815] = 3'b110;
        rom_memory[50816] = 3'b110;
        rom_memory[50817] = 3'b110;
        rom_memory[50818] = 3'b110;
        rom_memory[50819] = 3'b110;
        rom_memory[50820] = 3'b110;
        rom_memory[50821] = 3'b110;
        rom_memory[50822] = 3'b110;
        rom_memory[50823] = 3'b110;
        rom_memory[50824] = 3'b110;
        rom_memory[50825] = 3'b110;
        rom_memory[50826] = 3'b110;
        rom_memory[50827] = 3'b110;
        rom_memory[50828] = 3'b110;
        rom_memory[50829] = 3'b110;
        rom_memory[50830] = 3'b110;
        rom_memory[50831] = 3'b110;
        rom_memory[50832] = 3'b110;
        rom_memory[50833] = 3'b110;
        rom_memory[50834] = 3'b110;
        rom_memory[50835] = 3'b110;
        rom_memory[50836] = 3'b110;
        rom_memory[50837] = 3'b110;
        rom_memory[50838] = 3'b110;
        rom_memory[50839] = 3'b110;
        rom_memory[50840] = 3'b110;
        rom_memory[50841] = 3'b110;
        rom_memory[50842] = 3'b110;
        rom_memory[50843] = 3'b110;
        rom_memory[50844] = 3'b110;
        rom_memory[50845] = 3'b110;
        rom_memory[50846] = 3'b110;
        rom_memory[50847] = 3'b110;
        rom_memory[50848] = 3'b110;
        rom_memory[50849] = 3'b110;
        rom_memory[50850] = 3'b110;
        rom_memory[50851] = 3'b110;
        rom_memory[50852] = 3'b110;
        rom_memory[50853] = 3'b110;
        rom_memory[50854] = 3'b110;
        rom_memory[50855] = 3'b110;
        rom_memory[50856] = 3'b110;
        rom_memory[50857] = 3'b110;
        rom_memory[50858] = 3'b110;
        rom_memory[50859] = 3'b110;
        rom_memory[50860] = 3'b110;
        rom_memory[50861] = 3'b110;
        rom_memory[50862] = 3'b110;
        rom_memory[50863] = 3'b110;
        rom_memory[50864] = 3'b110;
        rom_memory[50865] = 3'b110;
        rom_memory[50866] = 3'b110;
        rom_memory[50867] = 3'b110;
        rom_memory[50868] = 3'b110;
        rom_memory[50869] = 3'b110;
        rom_memory[50870] = 3'b110;
        rom_memory[50871] = 3'b110;
        rom_memory[50872] = 3'b110;
        rom_memory[50873] = 3'b110;
        rom_memory[50874] = 3'b110;
        rom_memory[50875] = 3'b110;
        rom_memory[50876] = 3'b110;
        rom_memory[50877] = 3'b110;
        rom_memory[50878] = 3'b110;
        rom_memory[50879] = 3'b110;
        rom_memory[50880] = 3'b110;
        rom_memory[50881] = 3'b110;
        rom_memory[50882] = 3'b110;
        rom_memory[50883] = 3'b110;
        rom_memory[50884] = 3'b110;
        rom_memory[50885] = 3'b110;
        rom_memory[50886] = 3'b110;
        rom_memory[50887] = 3'b110;
        rom_memory[50888] = 3'b110;
        rom_memory[50889] = 3'b110;
        rom_memory[50890] = 3'b111;
        rom_memory[50891] = 3'b111;
        rom_memory[50892] = 3'b110;
        rom_memory[50893] = 3'b110;
        rom_memory[50894] = 3'b110;
        rom_memory[50895] = 3'b110;
        rom_memory[50896] = 3'b110;
        rom_memory[50897] = 3'b110;
        rom_memory[50898] = 3'b100;
        rom_memory[50899] = 3'b100;
        rom_memory[50900] = 3'b100;
        rom_memory[50901] = 3'b100;
        rom_memory[50902] = 3'b100;
        rom_memory[50903] = 3'b100;
        rom_memory[50904] = 3'b100;
        rom_memory[50905] = 3'b100;
        rom_memory[50906] = 3'b100;
        rom_memory[50907] = 3'b110;
        rom_memory[50908] = 3'b110;
        rom_memory[50909] = 3'b110;
        rom_memory[50910] = 3'b110;
        rom_memory[50911] = 3'b110;
        rom_memory[50912] = 3'b110;
        rom_memory[50913] = 3'b110;
        rom_memory[50914] = 3'b110;
        rom_memory[50915] = 3'b110;
        rom_memory[50916] = 3'b110;
        rom_memory[50917] = 3'b110;
        rom_memory[50918] = 3'b110;
        rom_memory[50919] = 3'b110;
        rom_memory[50920] = 3'b110;
        rom_memory[50921] = 3'b110;
        rom_memory[50922] = 3'b110;
        rom_memory[50923] = 3'b110;
        rom_memory[50924] = 3'b110;
        rom_memory[50925] = 3'b111;
        rom_memory[50926] = 3'b111;
        rom_memory[50927] = 3'b111;
        rom_memory[50928] = 3'b110;
        rom_memory[50929] = 3'b100;
        rom_memory[50930] = 3'b100;
        rom_memory[50931] = 3'b000;
        rom_memory[50932] = 3'b000;
        rom_memory[50933] = 3'b100;
        rom_memory[50934] = 3'b110;
        rom_memory[50935] = 3'b111;
        rom_memory[50936] = 3'b111;
        rom_memory[50937] = 3'b111;
        rom_memory[50938] = 3'b111;
        rom_memory[50939] = 3'b111;
        rom_memory[50940] = 3'b111;
        rom_memory[50941] = 3'b111;
        rom_memory[50942] = 3'b111;
        rom_memory[50943] = 3'b111;
        rom_memory[50944] = 3'b111;
        rom_memory[50945] = 3'b111;
        rom_memory[50946] = 3'b000;
        rom_memory[50947] = 3'b111;
        rom_memory[50948] = 3'b111;
        rom_memory[50949] = 3'b111;
        rom_memory[50950] = 3'b111;
        rom_memory[50951] = 3'b111;
        rom_memory[50952] = 3'b111;
        rom_memory[50953] = 3'b110;
        rom_memory[50954] = 3'b100;
        rom_memory[50955] = 3'b000;
        rom_memory[50956] = 3'b000;
        rom_memory[50957] = 3'b000;
        rom_memory[50958] = 3'b000;
        rom_memory[50959] = 3'b000;
        rom_memory[50960] = 3'b000;
        rom_memory[50961] = 3'b000;
        rom_memory[50962] = 3'b000;
        rom_memory[50963] = 3'b000;
        rom_memory[50964] = 3'b000;
        rom_memory[50965] = 3'b111;
        rom_memory[50966] = 3'b111;
        rom_memory[50967] = 3'b111;
        rom_memory[50968] = 3'b111;
        rom_memory[50969] = 3'b110;
        rom_memory[50970] = 3'b111;
        rom_memory[50971] = 3'b111;
        rom_memory[50972] = 3'b111;
        rom_memory[50973] = 3'b111;
        rom_memory[50974] = 3'b111;
        rom_memory[50975] = 3'b000;
        rom_memory[50976] = 3'b000;
        rom_memory[50977] = 3'b100;
        rom_memory[50978] = 3'b100;
        rom_memory[50979] = 3'b100;
        rom_memory[50980] = 3'b110;
        rom_memory[50981] = 3'b111;
        rom_memory[50982] = 3'b111;
        rom_memory[50983] = 3'b111;
        rom_memory[50984] = 3'b111;
        rom_memory[50985] = 3'b111;
        rom_memory[50986] = 3'b111;
        rom_memory[50987] = 3'b101;
        rom_memory[50988] = 3'b101;
        rom_memory[50989] = 3'b100;
        rom_memory[50990] = 3'b100;
        rom_memory[50991] = 3'b000;
        rom_memory[50992] = 3'b000;
        rom_memory[50993] = 3'b000;
        rom_memory[50994] = 3'b000;
        rom_memory[50995] = 3'b000;
        rom_memory[50996] = 3'b100;
        rom_memory[50997] = 3'b100;
        rom_memory[50998] = 3'b111;
        rom_memory[50999] = 3'b111;
        rom_memory[51000] = 3'b111;
        rom_memory[51001] = 3'b111;
        rom_memory[51002] = 3'b111;
        rom_memory[51003] = 3'b111;
        rom_memory[51004] = 3'b111;
        rom_memory[51005] = 3'b110;
        rom_memory[51006] = 3'b110;
        rom_memory[51007] = 3'b110;
        rom_memory[51008] = 3'b110;
        rom_memory[51009] = 3'b110;
        rom_memory[51010] = 3'b110;
        rom_memory[51011] = 3'b110;
        rom_memory[51012] = 3'b110;
        rom_memory[51013] = 3'b110;
        rom_memory[51014] = 3'b110;
        rom_memory[51015] = 3'b110;
        rom_memory[51016] = 3'b110;
        rom_memory[51017] = 3'b110;
        rom_memory[51018] = 3'b110;
        rom_memory[51019] = 3'b110;
        rom_memory[51020] = 3'b110;
        rom_memory[51021] = 3'b110;
        rom_memory[51022] = 3'b110;
        rom_memory[51023] = 3'b110;
        rom_memory[51024] = 3'b110;
        rom_memory[51025] = 3'b110;
        rom_memory[51026] = 3'b110;
        rom_memory[51027] = 3'b110;
        rom_memory[51028] = 3'b110;
        rom_memory[51029] = 3'b110;
        rom_memory[51030] = 3'b110;
        rom_memory[51031] = 3'b110;
        rom_memory[51032] = 3'b110;
        rom_memory[51033] = 3'b110;
        rom_memory[51034] = 3'b110;
        rom_memory[51035] = 3'b110;
        rom_memory[51036] = 3'b110;
        rom_memory[51037] = 3'b110;
        rom_memory[51038] = 3'b110;
        rom_memory[51039] = 3'b110;
        rom_memory[51040] = 3'b110;
        rom_memory[51041] = 3'b110;
        rom_memory[51042] = 3'b110;
        rom_memory[51043] = 3'b110;
        rom_memory[51044] = 3'b110;
        rom_memory[51045] = 3'b110;
        rom_memory[51046] = 3'b110;
        rom_memory[51047] = 3'b110;
        rom_memory[51048] = 3'b110;
        rom_memory[51049] = 3'b110;
        rom_memory[51050] = 3'b110;
        rom_memory[51051] = 3'b110;
        rom_memory[51052] = 3'b110;
        rom_memory[51053] = 3'b110;
        rom_memory[51054] = 3'b110;
        rom_memory[51055] = 3'b110;
        rom_memory[51056] = 3'b110;
        rom_memory[51057] = 3'b110;
        rom_memory[51058] = 3'b110;
        rom_memory[51059] = 3'b110;
        rom_memory[51060] = 3'b110;
        rom_memory[51061] = 3'b110;
        rom_memory[51062] = 3'b110;
        rom_memory[51063] = 3'b110;
        rom_memory[51064] = 3'b110;
        rom_memory[51065] = 3'b110;
        rom_memory[51066] = 3'b110;
        rom_memory[51067] = 3'b110;
        rom_memory[51068] = 3'b110;
        rom_memory[51069] = 3'b110;
        rom_memory[51070] = 3'b110;
        rom_memory[51071] = 3'b110;
        rom_memory[51072] = 3'b110;
        rom_memory[51073] = 3'b110;
        rom_memory[51074] = 3'b110;
        rom_memory[51075] = 3'b110;
        rom_memory[51076] = 3'b110;
        rom_memory[51077] = 3'b110;
        rom_memory[51078] = 3'b110;
        rom_memory[51079] = 3'b110;
        rom_memory[51080] = 3'b110;
        rom_memory[51081] = 3'b110;
        rom_memory[51082] = 3'b110;
        rom_memory[51083] = 3'b110;
        rom_memory[51084] = 3'b110;
        rom_memory[51085] = 3'b110;
        rom_memory[51086] = 3'b110;
        rom_memory[51087] = 3'b110;
        rom_memory[51088] = 3'b110;
        rom_memory[51089] = 3'b110;
        rom_memory[51090] = 3'b110;
        rom_memory[51091] = 3'b110;
        rom_memory[51092] = 3'b110;
        rom_memory[51093] = 3'b110;
        rom_memory[51094] = 3'b110;
        rom_memory[51095] = 3'b110;
        rom_memory[51096] = 3'b110;
        rom_memory[51097] = 3'b110;
        rom_memory[51098] = 3'b110;
        rom_memory[51099] = 3'b110;
        rom_memory[51100] = 3'b110;
        rom_memory[51101] = 3'b110;
        rom_memory[51102] = 3'b110;
        rom_memory[51103] = 3'b110;
        rom_memory[51104] = 3'b110;
        rom_memory[51105] = 3'b110;
        rom_memory[51106] = 3'b110;
        rom_memory[51107] = 3'b110;
        rom_memory[51108] = 3'b110;
        rom_memory[51109] = 3'b110;
        rom_memory[51110] = 3'b110;
        rom_memory[51111] = 3'b110;
        rom_memory[51112] = 3'b110;
        rom_memory[51113] = 3'b110;
        rom_memory[51114] = 3'b110;
        rom_memory[51115] = 3'b110;
        rom_memory[51116] = 3'b110;
        rom_memory[51117] = 3'b110;
        rom_memory[51118] = 3'b110;
        rom_memory[51119] = 3'b110;
        rom_memory[51120] = 3'b110;
        rom_memory[51121] = 3'b110;
        rom_memory[51122] = 3'b110;
        rom_memory[51123] = 3'b110;
        rom_memory[51124] = 3'b110;
        rom_memory[51125] = 3'b110;
        rom_memory[51126] = 3'b110;
        rom_memory[51127] = 3'b110;
        rom_memory[51128] = 3'b110;
        rom_memory[51129] = 3'b110;
        rom_memory[51130] = 3'b111;
        rom_memory[51131] = 3'b111;
        rom_memory[51132] = 3'b110;
        rom_memory[51133] = 3'b110;
        rom_memory[51134] = 3'b110;
        rom_memory[51135] = 3'b110;
        rom_memory[51136] = 3'b110;
        rom_memory[51137] = 3'b110;
        rom_memory[51138] = 3'b100;
        rom_memory[51139] = 3'b100;
        rom_memory[51140] = 3'b100;
        rom_memory[51141] = 3'b100;
        rom_memory[51142] = 3'b100;
        rom_memory[51143] = 3'b100;
        rom_memory[51144] = 3'b100;
        rom_memory[51145] = 3'b100;
        rom_memory[51146] = 3'b100;
        rom_memory[51147] = 3'b100;
        rom_memory[51148] = 3'b110;
        rom_memory[51149] = 3'b110;
        rom_memory[51150] = 3'b110;
        rom_memory[51151] = 3'b110;
        rom_memory[51152] = 3'b110;
        rom_memory[51153] = 3'b110;
        rom_memory[51154] = 3'b110;
        rom_memory[51155] = 3'b110;
        rom_memory[51156] = 3'b110;
        rom_memory[51157] = 3'b110;
        rom_memory[51158] = 3'b110;
        rom_memory[51159] = 3'b110;
        rom_memory[51160] = 3'b110;
        rom_memory[51161] = 3'b110;
        rom_memory[51162] = 3'b110;
        rom_memory[51163] = 3'b110;
        rom_memory[51164] = 3'b111;
        rom_memory[51165] = 3'b111;
        rom_memory[51166] = 3'b111;
        rom_memory[51167] = 3'b111;
        rom_memory[51168] = 3'b110;
        rom_memory[51169] = 3'b100;
        rom_memory[51170] = 3'b000;
        rom_memory[51171] = 3'b000;
        rom_memory[51172] = 3'b000;
        rom_memory[51173] = 3'b100;
        rom_memory[51174] = 3'b110;
        rom_memory[51175] = 3'b111;
        rom_memory[51176] = 3'b111;
        rom_memory[51177] = 3'b111;
        rom_memory[51178] = 3'b111;
        rom_memory[51179] = 3'b111;
        rom_memory[51180] = 3'b111;
        rom_memory[51181] = 3'b111;
        rom_memory[51182] = 3'b110;
        rom_memory[51183] = 3'b111;
        rom_memory[51184] = 3'b110;
        rom_memory[51185] = 3'b111;
        rom_memory[51186] = 3'b000;
        rom_memory[51187] = 3'b100;
        rom_memory[51188] = 3'b100;
        rom_memory[51189] = 3'b111;
        rom_memory[51190] = 3'b110;
        rom_memory[51191] = 3'b110;
        rom_memory[51192] = 3'b111;
        rom_memory[51193] = 3'b100;
        rom_memory[51194] = 3'b000;
        rom_memory[51195] = 3'b000;
        rom_memory[51196] = 3'b000;
        rom_memory[51197] = 3'b000;
        rom_memory[51198] = 3'b000;
        rom_memory[51199] = 3'b000;
        rom_memory[51200] = 3'b000;
        rom_memory[51201] = 3'b000;
        rom_memory[51202] = 3'b000;
        rom_memory[51203] = 3'b000;
        rom_memory[51204] = 3'b100;
        rom_memory[51205] = 3'b111;
        rom_memory[51206] = 3'b111;
        rom_memory[51207] = 3'b111;
        rom_memory[51208] = 3'b111;
        rom_memory[51209] = 3'b110;
        rom_memory[51210] = 3'b110;
        rom_memory[51211] = 3'b111;
        rom_memory[51212] = 3'b111;
        rom_memory[51213] = 3'b111;
        rom_memory[51214] = 3'b111;
        rom_memory[51215] = 3'b100;
        rom_memory[51216] = 3'b110;
        rom_memory[51217] = 3'b110;
        rom_memory[51218] = 3'b111;
        rom_memory[51219] = 3'b110;
        rom_memory[51220] = 3'b110;
        rom_memory[51221] = 3'b110;
        rom_memory[51222] = 3'b110;
        rom_memory[51223] = 3'b111;
        rom_memory[51224] = 3'b111;
        rom_memory[51225] = 3'b111;
        rom_memory[51226] = 3'b111;
        rom_memory[51227] = 3'b111;
        rom_memory[51228] = 3'b111;
        rom_memory[51229] = 3'b100;
        rom_memory[51230] = 3'b100;
        rom_memory[51231] = 3'b100;
        rom_memory[51232] = 3'b000;
        rom_memory[51233] = 3'b000;
        rom_memory[51234] = 3'b000;
        rom_memory[51235] = 3'b000;
        rom_memory[51236] = 3'b000;
        rom_memory[51237] = 3'b100;
        rom_memory[51238] = 3'b111;
        rom_memory[51239] = 3'b111;
        rom_memory[51240] = 3'b111;
        rom_memory[51241] = 3'b111;
        rom_memory[51242] = 3'b111;
        rom_memory[51243] = 3'b111;
        rom_memory[51244] = 3'b111;
        rom_memory[51245] = 3'b110;
        rom_memory[51246] = 3'b110;
        rom_memory[51247] = 3'b110;
        rom_memory[51248] = 3'b110;
        rom_memory[51249] = 3'b110;
        rom_memory[51250] = 3'b110;
        rom_memory[51251] = 3'b110;
        rom_memory[51252] = 3'b110;
        rom_memory[51253] = 3'b110;
        rom_memory[51254] = 3'b110;
        rom_memory[51255] = 3'b110;
        rom_memory[51256] = 3'b110;
        rom_memory[51257] = 3'b110;
        rom_memory[51258] = 3'b110;
        rom_memory[51259] = 3'b110;
        rom_memory[51260] = 3'b110;
        rom_memory[51261] = 3'b110;
        rom_memory[51262] = 3'b110;
        rom_memory[51263] = 3'b110;
        rom_memory[51264] = 3'b110;
        rom_memory[51265] = 3'b110;
        rom_memory[51266] = 3'b110;
        rom_memory[51267] = 3'b110;
        rom_memory[51268] = 3'b110;
        rom_memory[51269] = 3'b110;
        rom_memory[51270] = 3'b110;
        rom_memory[51271] = 3'b110;
        rom_memory[51272] = 3'b110;
        rom_memory[51273] = 3'b110;
        rom_memory[51274] = 3'b110;
        rom_memory[51275] = 3'b110;
        rom_memory[51276] = 3'b110;
        rom_memory[51277] = 3'b110;
        rom_memory[51278] = 3'b110;
        rom_memory[51279] = 3'b110;
        rom_memory[51280] = 3'b110;
        rom_memory[51281] = 3'b110;
        rom_memory[51282] = 3'b110;
        rom_memory[51283] = 3'b110;
        rom_memory[51284] = 3'b110;
        rom_memory[51285] = 3'b110;
        rom_memory[51286] = 3'b110;
        rom_memory[51287] = 3'b111;
        rom_memory[51288] = 3'b111;
        rom_memory[51289] = 3'b111;
        rom_memory[51290] = 3'b111;
        rom_memory[51291] = 3'b111;
        rom_memory[51292] = 3'b111;
        rom_memory[51293] = 3'b111;
        rom_memory[51294] = 3'b110;
        rom_memory[51295] = 3'b111;
        rom_memory[51296] = 3'b111;
        rom_memory[51297] = 3'b111;
        rom_memory[51298] = 3'b110;
        rom_memory[51299] = 3'b110;
        rom_memory[51300] = 3'b110;
        rom_memory[51301] = 3'b111;
        rom_memory[51302] = 3'b110;
        rom_memory[51303] = 3'b110;
        rom_memory[51304] = 3'b110;
        rom_memory[51305] = 3'b110;
        rom_memory[51306] = 3'b110;
        rom_memory[51307] = 3'b110;
        rom_memory[51308] = 3'b110;
        rom_memory[51309] = 3'b110;
        rom_memory[51310] = 3'b110;
        rom_memory[51311] = 3'b110;
        rom_memory[51312] = 3'b110;
        rom_memory[51313] = 3'b110;
        rom_memory[51314] = 3'b110;
        rom_memory[51315] = 3'b110;
        rom_memory[51316] = 3'b110;
        rom_memory[51317] = 3'b110;
        rom_memory[51318] = 3'b110;
        rom_memory[51319] = 3'b110;
        rom_memory[51320] = 3'b110;
        rom_memory[51321] = 3'b110;
        rom_memory[51322] = 3'b110;
        rom_memory[51323] = 3'b110;
        rom_memory[51324] = 3'b110;
        rom_memory[51325] = 3'b110;
        rom_memory[51326] = 3'b110;
        rom_memory[51327] = 3'b110;
        rom_memory[51328] = 3'b110;
        rom_memory[51329] = 3'b110;
        rom_memory[51330] = 3'b110;
        rom_memory[51331] = 3'b110;
        rom_memory[51332] = 3'b110;
        rom_memory[51333] = 3'b110;
        rom_memory[51334] = 3'b110;
        rom_memory[51335] = 3'b110;
        rom_memory[51336] = 3'b110;
        rom_memory[51337] = 3'b110;
        rom_memory[51338] = 3'b111;
        rom_memory[51339] = 3'b110;
        rom_memory[51340] = 3'b110;
        rom_memory[51341] = 3'b110;
        rom_memory[51342] = 3'b110;
        rom_memory[51343] = 3'b110;
        rom_memory[51344] = 3'b110;
        rom_memory[51345] = 3'b110;
        rom_memory[51346] = 3'b110;
        rom_memory[51347] = 3'b110;
        rom_memory[51348] = 3'b110;
        rom_memory[51349] = 3'b110;
        rom_memory[51350] = 3'b110;
        rom_memory[51351] = 3'b110;
        rom_memory[51352] = 3'b110;
        rom_memory[51353] = 3'b110;
        rom_memory[51354] = 3'b110;
        rom_memory[51355] = 3'b110;
        rom_memory[51356] = 3'b110;
        rom_memory[51357] = 3'b110;
        rom_memory[51358] = 3'b111;
        rom_memory[51359] = 3'b110;
        rom_memory[51360] = 3'b110;
        rom_memory[51361] = 3'b110;
        rom_memory[51362] = 3'b110;
        rom_memory[51363] = 3'b110;
        rom_memory[51364] = 3'b110;
        rom_memory[51365] = 3'b110;
        rom_memory[51366] = 3'b110;
        rom_memory[51367] = 3'b110;
        rom_memory[51368] = 3'b110;
        rom_memory[51369] = 3'b110;
        rom_memory[51370] = 3'b111;
        rom_memory[51371] = 3'b111;
        rom_memory[51372] = 3'b110;
        rom_memory[51373] = 3'b110;
        rom_memory[51374] = 3'b110;
        rom_memory[51375] = 3'b110;
        rom_memory[51376] = 3'b110;
        rom_memory[51377] = 3'b110;
        rom_memory[51378] = 3'b100;
        rom_memory[51379] = 3'b100;
        rom_memory[51380] = 3'b100;
        rom_memory[51381] = 3'b100;
        rom_memory[51382] = 3'b100;
        rom_memory[51383] = 3'b100;
        rom_memory[51384] = 3'b100;
        rom_memory[51385] = 3'b100;
        rom_memory[51386] = 3'b100;
        rom_memory[51387] = 3'b100;
        rom_memory[51388] = 3'b100;
        rom_memory[51389] = 3'b110;
        rom_memory[51390] = 3'b110;
        rom_memory[51391] = 3'b110;
        rom_memory[51392] = 3'b110;
        rom_memory[51393] = 3'b110;
        rom_memory[51394] = 3'b110;
        rom_memory[51395] = 3'b110;
        rom_memory[51396] = 3'b110;
        rom_memory[51397] = 3'b110;
        rom_memory[51398] = 3'b110;
        rom_memory[51399] = 3'b111;
        rom_memory[51400] = 3'b110;
        rom_memory[51401] = 3'b110;
        rom_memory[51402] = 3'b110;
        rom_memory[51403] = 3'b110;
        rom_memory[51404] = 3'b110;
        rom_memory[51405] = 3'b110;
        rom_memory[51406] = 3'b111;
        rom_memory[51407] = 3'b111;
        rom_memory[51408] = 3'b110;
        rom_memory[51409] = 3'b000;
        rom_memory[51410] = 3'b000;
        rom_memory[51411] = 3'b000;
        rom_memory[51412] = 3'b000;
        rom_memory[51413] = 3'b110;
        rom_memory[51414] = 3'b111;
        rom_memory[51415] = 3'b111;
        rom_memory[51416] = 3'b111;
        rom_memory[51417] = 3'b111;
        rom_memory[51418] = 3'b111;
        rom_memory[51419] = 3'b111;
        rom_memory[51420] = 3'b111;
        rom_memory[51421] = 3'b110;
        rom_memory[51422] = 3'b110;
        rom_memory[51423] = 3'b111;
        rom_memory[51424] = 3'b110;
        rom_memory[51425] = 3'b100;
        rom_memory[51426] = 3'b000;
        rom_memory[51427] = 3'b100;
        rom_memory[51428] = 3'b100;
        rom_memory[51429] = 3'b100;
        rom_memory[51430] = 3'b100;
        rom_memory[51431] = 3'b100;
        rom_memory[51432] = 3'b110;
        rom_memory[51433] = 3'b110;
        rom_memory[51434] = 3'b100;
        rom_memory[51435] = 3'b000;
        rom_memory[51436] = 3'b000;
        rom_memory[51437] = 3'b000;
        rom_memory[51438] = 3'b000;
        rom_memory[51439] = 3'b000;
        rom_memory[51440] = 3'b000;
        rom_memory[51441] = 3'b000;
        rom_memory[51442] = 3'b000;
        rom_memory[51443] = 3'b000;
        rom_memory[51444] = 3'b110;
        rom_memory[51445] = 3'b111;
        rom_memory[51446] = 3'b111;
        rom_memory[51447] = 3'b111;
        rom_memory[51448] = 3'b111;
        rom_memory[51449] = 3'b111;
        rom_memory[51450] = 3'b111;
        rom_memory[51451] = 3'b111;
        rom_memory[51452] = 3'b111;
        rom_memory[51453] = 3'b111;
        rom_memory[51454] = 3'b111;
        rom_memory[51455] = 3'b111;
        rom_memory[51456] = 3'b111;
        rom_memory[51457] = 3'b111;
        rom_memory[51458] = 3'b111;
        rom_memory[51459] = 3'b111;
        rom_memory[51460] = 3'b111;
        rom_memory[51461] = 3'b111;
        rom_memory[51462] = 3'b111;
        rom_memory[51463] = 3'b110;
        rom_memory[51464] = 3'b110;
        rom_memory[51465] = 3'b111;
        rom_memory[51466] = 3'b101;
        rom_memory[51467] = 3'b111;
        rom_memory[51468] = 3'b111;
        rom_memory[51469] = 3'b100;
        rom_memory[51470] = 3'b100;
        rom_memory[51471] = 3'b100;
        rom_memory[51472] = 3'b000;
        rom_memory[51473] = 3'b000;
        rom_memory[51474] = 3'b000;
        rom_memory[51475] = 3'b000;
        rom_memory[51476] = 3'b000;
        rom_memory[51477] = 3'b100;
        rom_memory[51478] = 3'b100;
        rom_memory[51479] = 3'b111;
        rom_memory[51480] = 3'b111;
        rom_memory[51481] = 3'b111;
        rom_memory[51482] = 3'b111;
        rom_memory[51483] = 3'b111;
        rom_memory[51484] = 3'b111;
        rom_memory[51485] = 3'b110;
        rom_memory[51486] = 3'b110;
        rom_memory[51487] = 3'b110;
        rom_memory[51488] = 3'b110;
        rom_memory[51489] = 3'b110;
        rom_memory[51490] = 3'b110;
        rom_memory[51491] = 3'b110;
        rom_memory[51492] = 3'b110;
        rom_memory[51493] = 3'b110;
        rom_memory[51494] = 3'b110;
        rom_memory[51495] = 3'b110;
        rom_memory[51496] = 3'b110;
        rom_memory[51497] = 3'b110;
        rom_memory[51498] = 3'b110;
        rom_memory[51499] = 3'b110;
        rom_memory[51500] = 3'b110;
        rom_memory[51501] = 3'b110;
        rom_memory[51502] = 3'b110;
        rom_memory[51503] = 3'b110;
        rom_memory[51504] = 3'b110;
        rom_memory[51505] = 3'b110;
        rom_memory[51506] = 3'b110;
        rom_memory[51507] = 3'b110;
        rom_memory[51508] = 3'b110;
        rom_memory[51509] = 3'b110;
        rom_memory[51510] = 3'b110;
        rom_memory[51511] = 3'b110;
        rom_memory[51512] = 3'b110;
        rom_memory[51513] = 3'b110;
        rom_memory[51514] = 3'b110;
        rom_memory[51515] = 3'b110;
        rom_memory[51516] = 3'b110;
        rom_memory[51517] = 3'b110;
        rom_memory[51518] = 3'b110;
        rom_memory[51519] = 3'b110;
        rom_memory[51520] = 3'b111;
        rom_memory[51521] = 3'b111;
        rom_memory[51522] = 3'b111;
        rom_memory[51523] = 3'b111;
        rom_memory[51524] = 3'b111;
        rom_memory[51525] = 3'b111;
        rom_memory[51526] = 3'b111;
        rom_memory[51527] = 3'b111;
        rom_memory[51528] = 3'b111;
        rom_memory[51529] = 3'b111;
        rom_memory[51530] = 3'b111;
        rom_memory[51531] = 3'b111;
        rom_memory[51532] = 3'b111;
        rom_memory[51533] = 3'b111;
        rom_memory[51534] = 3'b111;
        rom_memory[51535] = 3'b111;
        rom_memory[51536] = 3'b111;
        rom_memory[51537] = 3'b111;
        rom_memory[51538] = 3'b111;
        rom_memory[51539] = 3'b111;
        rom_memory[51540] = 3'b111;
        rom_memory[51541] = 3'b111;
        rom_memory[51542] = 3'b111;
        rom_memory[51543] = 3'b111;
        rom_memory[51544] = 3'b111;
        rom_memory[51545] = 3'b111;
        rom_memory[51546] = 3'b111;
        rom_memory[51547] = 3'b111;
        rom_memory[51548] = 3'b111;
        rom_memory[51549] = 3'b111;
        rom_memory[51550] = 3'b111;
        rom_memory[51551] = 3'b111;
        rom_memory[51552] = 3'b111;
        rom_memory[51553] = 3'b111;
        rom_memory[51554] = 3'b111;
        rom_memory[51555] = 3'b111;
        rom_memory[51556] = 3'b111;
        rom_memory[51557] = 3'b111;
        rom_memory[51558] = 3'b111;
        rom_memory[51559] = 3'b111;
        rom_memory[51560] = 3'b111;
        rom_memory[51561] = 3'b111;
        rom_memory[51562] = 3'b111;
        rom_memory[51563] = 3'b111;
        rom_memory[51564] = 3'b111;
        rom_memory[51565] = 3'b111;
        rom_memory[51566] = 3'b111;
        rom_memory[51567] = 3'b111;
        rom_memory[51568] = 3'b111;
        rom_memory[51569] = 3'b111;
        rom_memory[51570] = 3'b111;
        rom_memory[51571] = 3'b111;
        rom_memory[51572] = 3'b111;
        rom_memory[51573] = 3'b111;
        rom_memory[51574] = 3'b111;
        rom_memory[51575] = 3'b111;
        rom_memory[51576] = 3'b111;
        rom_memory[51577] = 3'b111;
        rom_memory[51578] = 3'b111;
        rom_memory[51579] = 3'b111;
        rom_memory[51580] = 3'b111;
        rom_memory[51581] = 3'b111;
        rom_memory[51582] = 3'b111;
        rom_memory[51583] = 3'b111;
        rom_memory[51584] = 3'b111;
        rom_memory[51585] = 3'b111;
        rom_memory[51586] = 3'b111;
        rom_memory[51587] = 3'b111;
        rom_memory[51588] = 3'b111;
        rom_memory[51589] = 3'b111;
        rom_memory[51590] = 3'b111;
        rom_memory[51591] = 3'b111;
        rom_memory[51592] = 3'b111;
        rom_memory[51593] = 3'b111;
        rom_memory[51594] = 3'b111;
        rom_memory[51595] = 3'b111;
        rom_memory[51596] = 3'b111;
        rom_memory[51597] = 3'b111;
        rom_memory[51598] = 3'b111;
        rom_memory[51599] = 3'b111;
        rom_memory[51600] = 3'b110;
        rom_memory[51601] = 3'b110;
        rom_memory[51602] = 3'b110;
        rom_memory[51603] = 3'b110;
        rom_memory[51604] = 3'b110;
        rom_memory[51605] = 3'b110;
        rom_memory[51606] = 3'b110;
        rom_memory[51607] = 3'b110;
        rom_memory[51608] = 3'b111;
        rom_memory[51609] = 3'b111;
        rom_memory[51610] = 3'b111;
        rom_memory[51611] = 3'b111;
        rom_memory[51612] = 3'b110;
        rom_memory[51613] = 3'b110;
        rom_memory[51614] = 3'b110;
        rom_memory[51615] = 3'b110;
        rom_memory[51616] = 3'b110;
        rom_memory[51617] = 3'b110;
        rom_memory[51618] = 3'b100;
        rom_memory[51619] = 3'b100;
        rom_memory[51620] = 3'b100;
        rom_memory[51621] = 3'b100;
        rom_memory[51622] = 3'b100;
        rom_memory[51623] = 3'b100;
        rom_memory[51624] = 3'b100;
        rom_memory[51625] = 3'b100;
        rom_memory[51626] = 3'b100;
        rom_memory[51627] = 3'b100;
        rom_memory[51628] = 3'b100;
        rom_memory[51629] = 3'b100;
        rom_memory[51630] = 3'b110;
        rom_memory[51631] = 3'b110;
        rom_memory[51632] = 3'b110;
        rom_memory[51633] = 3'b110;
        rom_memory[51634] = 3'b110;
        rom_memory[51635] = 3'b110;
        rom_memory[51636] = 3'b110;
        rom_memory[51637] = 3'b110;
        rom_memory[51638] = 3'b110;
        rom_memory[51639] = 3'b111;
        rom_memory[51640] = 3'b111;
        rom_memory[51641] = 3'b111;
        rom_memory[51642] = 3'b110;
        rom_memory[51643] = 3'b110;
        rom_memory[51644] = 3'b110;
        rom_memory[51645] = 3'b110;
        rom_memory[51646] = 3'b111;
        rom_memory[51647] = 3'b111;
        rom_memory[51648] = 3'b111;
        rom_memory[51649] = 3'b100;
        rom_memory[51650] = 3'b100;
        rom_memory[51651] = 3'b100;
        rom_memory[51652] = 3'b000;
        rom_memory[51653] = 3'b110;
        rom_memory[51654] = 3'b111;
        rom_memory[51655] = 3'b111;
        rom_memory[51656] = 3'b111;
        rom_memory[51657] = 3'b111;
        rom_memory[51658] = 3'b111;
        rom_memory[51659] = 3'b111;
        rom_memory[51660] = 3'b111;
        rom_memory[51661] = 3'b110;
        rom_memory[51662] = 3'b110;
        rom_memory[51663] = 3'b110;
        rom_memory[51664] = 3'b110;
        rom_memory[51665] = 3'b000;
        rom_memory[51666] = 3'b000;
        rom_memory[51667] = 3'b100;
        rom_memory[51668] = 3'b111;
        rom_memory[51669] = 3'b100;
        rom_memory[51670] = 3'b100;
        rom_memory[51671] = 3'b110;
        rom_memory[51672] = 3'b111;
        rom_memory[51673] = 3'b110;
        rom_memory[51674] = 3'b110;
        rom_memory[51675] = 3'b100;
        rom_memory[51676] = 3'b100;
        rom_memory[51677] = 3'b100;
        rom_memory[51678] = 3'b100;
        rom_memory[51679] = 3'b000;
        rom_memory[51680] = 3'b000;
        rom_memory[51681] = 3'b000;
        rom_memory[51682] = 3'b000;
        rom_memory[51683] = 3'b100;
        rom_memory[51684] = 3'b110;
        rom_memory[51685] = 3'b111;
        rom_memory[51686] = 3'b111;
        rom_memory[51687] = 3'b111;
        rom_memory[51688] = 3'b111;
        rom_memory[51689] = 3'b111;
        rom_memory[51690] = 3'b111;
        rom_memory[51691] = 3'b111;
        rom_memory[51692] = 3'b111;
        rom_memory[51693] = 3'b111;
        rom_memory[51694] = 3'b111;
        rom_memory[51695] = 3'b111;
        rom_memory[51696] = 3'b111;
        rom_memory[51697] = 3'b111;
        rom_memory[51698] = 3'b111;
        rom_memory[51699] = 3'b111;
        rom_memory[51700] = 3'b111;
        rom_memory[51701] = 3'b111;
        rom_memory[51702] = 3'b111;
        rom_memory[51703] = 3'b111;
        rom_memory[51704] = 3'b110;
        rom_memory[51705] = 3'b110;
        rom_memory[51706] = 3'b111;
        rom_memory[51707] = 3'b111;
        rom_memory[51708] = 3'b100;
        rom_memory[51709] = 3'b100;
        rom_memory[51710] = 3'b100;
        rom_memory[51711] = 3'b100;
        rom_memory[51712] = 3'b100;
        rom_memory[51713] = 3'b000;
        rom_memory[51714] = 3'b000;
        rom_memory[51715] = 3'b000;
        rom_memory[51716] = 3'b000;
        rom_memory[51717] = 3'b000;
        rom_memory[51718] = 3'b100;
        rom_memory[51719] = 3'b111;
        rom_memory[51720] = 3'b111;
        rom_memory[51721] = 3'b111;
        rom_memory[51722] = 3'b111;
        rom_memory[51723] = 3'b111;
        rom_memory[51724] = 3'b111;
        rom_memory[51725] = 3'b111;
        rom_memory[51726] = 3'b110;
        rom_memory[51727] = 3'b110;
        rom_memory[51728] = 3'b110;
        rom_memory[51729] = 3'b110;
        rom_memory[51730] = 3'b110;
        rom_memory[51731] = 3'b110;
        rom_memory[51732] = 3'b110;
        rom_memory[51733] = 3'b110;
        rom_memory[51734] = 3'b110;
        rom_memory[51735] = 3'b110;
        rom_memory[51736] = 3'b110;
        rom_memory[51737] = 3'b110;
        rom_memory[51738] = 3'b110;
        rom_memory[51739] = 3'b110;
        rom_memory[51740] = 3'b110;
        rom_memory[51741] = 3'b110;
        rom_memory[51742] = 3'b110;
        rom_memory[51743] = 3'b110;
        rom_memory[51744] = 3'b110;
        rom_memory[51745] = 3'b110;
        rom_memory[51746] = 3'b110;
        rom_memory[51747] = 3'b110;
        rom_memory[51748] = 3'b110;
        rom_memory[51749] = 3'b110;
        rom_memory[51750] = 3'b110;
        rom_memory[51751] = 3'b110;
        rom_memory[51752] = 3'b110;
        rom_memory[51753] = 3'b110;
        rom_memory[51754] = 3'b110;
        rom_memory[51755] = 3'b110;
        rom_memory[51756] = 3'b110;
        rom_memory[51757] = 3'b110;
        rom_memory[51758] = 3'b110;
        rom_memory[51759] = 3'b111;
        rom_memory[51760] = 3'b111;
        rom_memory[51761] = 3'b111;
        rom_memory[51762] = 3'b111;
        rom_memory[51763] = 3'b111;
        rom_memory[51764] = 3'b111;
        rom_memory[51765] = 3'b111;
        rom_memory[51766] = 3'b111;
        rom_memory[51767] = 3'b111;
        rom_memory[51768] = 3'b111;
        rom_memory[51769] = 3'b111;
        rom_memory[51770] = 3'b111;
        rom_memory[51771] = 3'b111;
        rom_memory[51772] = 3'b111;
        rom_memory[51773] = 3'b111;
        rom_memory[51774] = 3'b111;
        rom_memory[51775] = 3'b111;
        rom_memory[51776] = 3'b111;
        rom_memory[51777] = 3'b111;
        rom_memory[51778] = 3'b111;
        rom_memory[51779] = 3'b111;
        rom_memory[51780] = 3'b111;
        rom_memory[51781] = 3'b111;
        rom_memory[51782] = 3'b111;
        rom_memory[51783] = 3'b111;
        rom_memory[51784] = 3'b111;
        rom_memory[51785] = 3'b111;
        rom_memory[51786] = 3'b111;
        rom_memory[51787] = 3'b111;
        rom_memory[51788] = 3'b111;
        rom_memory[51789] = 3'b111;
        rom_memory[51790] = 3'b111;
        rom_memory[51791] = 3'b111;
        rom_memory[51792] = 3'b111;
        rom_memory[51793] = 3'b111;
        rom_memory[51794] = 3'b111;
        rom_memory[51795] = 3'b111;
        rom_memory[51796] = 3'b111;
        rom_memory[51797] = 3'b111;
        rom_memory[51798] = 3'b111;
        rom_memory[51799] = 3'b111;
        rom_memory[51800] = 3'b111;
        rom_memory[51801] = 3'b111;
        rom_memory[51802] = 3'b111;
        rom_memory[51803] = 3'b111;
        rom_memory[51804] = 3'b111;
        rom_memory[51805] = 3'b111;
        rom_memory[51806] = 3'b111;
        rom_memory[51807] = 3'b111;
        rom_memory[51808] = 3'b111;
        rom_memory[51809] = 3'b111;
        rom_memory[51810] = 3'b111;
        rom_memory[51811] = 3'b111;
        rom_memory[51812] = 3'b111;
        rom_memory[51813] = 3'b111;
        rom_memory[51814] = 3'b111;
        rom_memory[51815] = 3'b111;
        rom_memory[51816] = 3'b111;
        rom_memory[51817] = 3'b111;
        rom_memory[51818] = 3'b111;
        rom_memory[51819] = 3'b111;
        rom_memory[51820] = 3'b111;
        rom_memory[51821] = 3'b111;
        rom_memory[51822] = 3'b111;
        rom_memory[51823] = 3'b111;
        rom_memory[51824] = 3'b111;
        rom_memory[51825] = 3'b111;
        rom_memory[51826] = 3'b111;
        rom_memory[51827] = 3'b111;
        rom_memory[51828] = 3'b111;
        rom_memory[51829] = 3'b111;
        rom_memory[51830] = 3'b111;
        rom_memory[51831] = 3'b111;
        rom_memory[51832] = 3'b111;
        rom_memory[51833] = 3'b111;
        rom_memory[51834] = 3'b111;
        rom_memory[51835] = 3'b111;
        rom_memory[51836] = 3'b111;
        rom_memory[51837] = 3'b111;
        rom_memory[51838] = 3'b111;
        rom_memory[51839] = 3'b111;
        rom_memory[51840] = 3'b110;
        rom_memory[51841] = 3'b110;
        rom_memory[51842] = 3'b110;
        rom_memory[51843] = 3'b110;
        rom_memory[51844] = 3'b110;
        rom_memory[51845] = 3'b110;
        rom_memory[51846] = 3'b110;
        rom_memory[51847] = 3'b110;
        rom_memory[51848] = 3'b111;
        rom_memory[51849] = 3'b111;
        rom_memory[51850] = 3'b111;
        rom_memory[51851] = 3'b111;
        rom_memory[51852] = 3'b110;
        rom_memory[51853] = 3'b110;
        rom_memory[51854] = 3'b110;
        rom_memory[51855] = 3'b110;
        rom_memory[51856] = 3'b110;
        rom_memory[51857] = 3'b110;
        rom_memory[51858] = 3'b100;
        rom_memory[51859] = 3'b100;
        rom_memory[51860] = 3'b100;
        rom_memory[51861] = 3'b100;
        rom_memory[51862] = 3'b100;
        rom_memory[51863] = 3'b100;
        rom_memory[51864] = 3'b100;
        rom_memory[51865] = 3'b100;
        rom_memory[51866] = 3'b100;
        rom_memory[51867] = 3'b100;
        rom_memory[51868] = 3'b100;
        rom_memory[51869] = 3'b100;
        rom_memory[51870] = 3'b110;
        rom_memory[51871] = 3'b110;
        rom_memory[51872] = 3'b110;
        rom_memory[51873] = 3'b110;
        rom_memory[51874] = 3'b110;
        rom_memory[51875] = 3'b110;
        rom_memory[51876] = 3'b111;
        rom_memory[51877] = 3'b111;
        rom_memory[51878] = 3'b111;
        rom_memory[51879] = 3'b111;
        rom_memory[51880] = 3'b111;
        rom_memory[51881] = 3'b111;
        rom_memory[51882] = 3'b111;
        rom_memory[51883] = 3'b110;
        rom_memory[51884] = 3'b110;
        rom_memory[51885] = 3'b110;
        rom_memory[51886] = 3'b111;
        rom_memory[51887] = 3'b111;
        rom_memory[51888] = 3'b111;
        rom_memory[51889] = 3'b111;
        rom_memory[51890] = 3'b000;
        rom_memory[51891] = 3'b000;
        rom_memory[51892] = 3'b000;
        rom_memory[51893] = 3'b100;
        rom_memory[51894] = 3'b111;
        rom_memory[51895] = 3'b111;
        rom_memory[51896] = 3'b111;
        rom_memory[51897] = 3'b111;
        rom_memory[51898] = 3'b111;
        rom_memory[51899] = 3'b111;
        rom_memory[51900] = 3'b111;
        rom_memory[51901] = 3'b110;
        rom_memory[51902] = 3'b110;
        rom_memory[51903] = 3'b110;
        rom_memory[51904] = 3'b110;
        rom_memory[51905] = 3'b000;
        rom_memory[51906] = 3'b000;
        rom_memory[51907] = 3'b000;
        rom_memory[51908] = 3'b111;
        rom_memory[51909] = 3'b110;
        rom_memory[51910] = 3'b100;
        rom_memory[51911] = 3'b111;
        rom_memory[51912] = 3'b110;
        rom_memory[51913] = 3'b110;
        rom_memory[51914] = 3'b110;
        rom_memory[51915] = 3'b100;
        rom_memory[51916] = 3'b100;
        rom_memory[51917] = 3'b100;
        rom_memory[51918] = 3'b100;
        rom_memory[51919] = 3'b100;
        rom_memory[51920] = 3'b100;
        rom_memory[51921] = 3'b000;
        rom_memory[51922] = 3'b100;
        rom_memory[51923] = 3'b110;
        rom_memory[51924] = 3'b111;
        rom_memory[51925] = 3'b111;
        rom_memory[51926] = 3'b111;
        rom_memory[51927] = 3'b111;
        rom_memory[51928] = 3'b111;
        rom_memory[51929] = 3'b111;
        rom_memory[51930] = 3'b111;
        rom_memory[51931] = 3'b111;
        rom_memory[51932] = 3'b111;
        rom_memory[51933] = 3'b111;
        rom_memory[51934] = 3'b111;
        rom_memory[51935] = 3'b111;
        rom_memory[51936] = 3'b111;
        rom_memory[51937] = 3'b111;
        rom_memory[51938] = 3'b111;
        rom_memory[51939] = 3'b111;
        rom_memory[51940] = 3'b111;
        rom_memory[51941] = 3'b110;
        rom_memory[51942] = 3'b110;
        rom_memory[51943] = 3'b111;
        rom_memory[51944] = 3'b111;
        rom_memory[51945] = 3'b111;
        rom_memory[51946] = 3'b111;
        rom_memory[51947] = 3'b111;
        rom_memory[51948] = 3'b100;
        rom_memory[51949] = 3'b100;
        rom_memory[51950] = 3'b100;
        rom_memory[51951] = 3'b100;
        rom_memory[51952] = 3'b100;
        rom_memory[51953] = 3'b100;
        rom_memory[51954] = 3'b000;
        rom_memory[51955] = 3'b000;
        rom_memory[51956] = 3'b000;
        rom_memory[51957] = 3'b000;
        rom_memory[51958] = 3'b100;
        rom_memory[51959] = 3'b100;
        rom_memory[51960] = 3'b111;
        rom_memory[51961] = 3'b111;
        rom_memory[51962] = 3'b111;
        rom_memory[51963] = 3'b111;
        rom_memory[51964] = 3'b111;
        rom_memory[51965] = 3'b111;
        rom_memory[51966] = 3'b110;
        rom_memory[51967] = 3'b110;
        rom_memory[51968] = 3'b110;
        rom_memory[51969] = 3'b110;
        rom_memory[51970] = 3'b110;
        rom_memory[51971] = 3'b110;
        rom_memory[51972] = 3'b110;
        rom_memory[51973] = 3'b110;
        rom_memory[51974] = 3'b110;
        rom_memory[51975] = 3'b110;
        rom_memory[51976] = 3'b110;
        rom_memory[51977] = 3'b110;
        rom_memory[51978] = 3'b110;
        rom_memory[51979] = 3'b110;
        rom_memory[51980] = 3'b110;
        rom_memory[51981] = 3'b110;
        rom_memory[51982] = 3'b110;
        rom_memory[51983] = 3'b110;
        rom_memory[51984] = 3'b110;
        rom_memory[51985] = 3'b110;
        rom_memory[51986] = 3'b110;
        rom_memory[51987] = 3'b110;
        rom_memory[51988] = 3'b110;
        rom_memory[51989] = 3'b110;
        rom_memory[51990] = 3'b110;
        rom_memory[51991] = 3'b110;
        rom_memory[51992] = 3'b110;
        rom_memory[51993] = 3'b110;
        rom_memory[51994] = 3'b110;
        rom_memory[51995] = 3'b110;
        rom_memory[51996] = 3'b110;
        rom_memory[51997] = 3'b110;
        rom_memory[51998] = 3'b110;
        rom_memory[51999] = 3'b111;
        rom_memory[52000] = 3'b111;
        rom_memory[52001] = 3'b111;
        rom_memory[52002] = 3'b111;
        rom_memory[52003] = 3'b111;
        rom_memory[52004] = 3'b111;
        rom_memory[52005] = 3'b111;
        rom_memory[52006] = 3'b111;
        rom_memory[52007] = 3'b111;
        rom_memory[52008] = 3'b111;
        rom_memory[52009] = 3'b111;
        rom_memory[52010] = 3'b111;
        rom_memory[52011] = 3'b111;
        rom_memory[52012] = 3'b111;
        rom_memory[52013] = 3'b111;
        rom_memory[52014] = 3'b111;
        rom_memory[52015] = 3'b111;
        rom_memory[52016] = 3'b111;
        rom_memory[52017] = 3'b111;
        rom_memory[52018] = 3'b111;
        rom_memory[52019] = 3'b111;
        rom_memory[52020] = 3'b111;
        rom_memory[52021] = 3'b111;
        rom_memory[52022] = 3'b111;
        rom_memory[52023] = 3'b111;
        rom_memory[52024] = 3'b111;
        rom_memory[52025] = 3'b111;
        rom_memory[52026] = 3'b111;
        rom_memory[52027] = 3'b111;
        rom_memory[52028] = 3'b111;
        rom_memory[52029] = 3'b111;
        rom_memory[52030] = 3'b111;
        rom_memory[52031] = 3'b111;
        rom_memory[52032] = 3'b111;
        rom_memory[52033] = 3'b111;
        rom_memory[52034] = 3'b111;
        rom_memory[52035] = 3'b111;
        rom_memory[52036] = 3'b111;
        rom_memory[52037] = 3'b111;
        rom_memory[52038] = 3'b111;
        rom_memory[52039] = 3'b111;
        rom_memory[52040] = 3'b111;
        rom_memory[52041] = 3'b111;
        rom_memory[52042] = 3'b111;
        rom_memory[52043] = 3'b111;
        rom_memory[52044] = 3'b111;
        rom_memory[52045] = 3'b111;
        rom_memory[52046] = 3'b111;
        rom_memory[52047] = 3'b111;
        rom_memory[52048] = 3'b111;
        rom_memory[52049] = 3'b111;
        rom_memory[52050] = 3'b111;
        rom_memory[52051] = 3'b111;
        rom_memory[52052] = 3'b111;
        rom_memory[52053] = 3'b111;
        rom_memory[52054] = 3'b111;
        rom_memory[52055] = 3'b111;
        rom_memory[52056] = 3'b111;
        rom_memory[52057] = 3'b111;
        rom_memory[52058] = 3'b111;
        rom_memory[52059] = 3'b111;
        rom_memory[52060] = 3'b111;
        rom_memory[52061] = 3'b111;
        rom_memory[52062] = 3'b111;
        rom_memory[52063] = 3'b111;
        rom_memory[52064] = 3'b111;
        rom_memory[52065] = 3'b111;
        rom_memory[52066] = 3'b111;
        rom_memory[52067] = 3'b111;
        rom_memory[52068] = 3'b111;
        rom_memory[52069] = 3'b111;
        rom_memory[52070] = 3'b111;
        rom_memory[52071] = 3'b111;
        rom_memory[52072] = 3'b111;
        rom_memory[52073] = 3'b111;
        rom_memory[52074] = 3'b111;
        rom_memory[52075] = 3'b111;
        rom_memory[52076] = 3'b111;
        rom_memory[52077] = 3'b111;
        rom_memory[52078] = 3'b111;
        rom_memory[52079] = 3'b111;
        rom_memory[52080] = 3'b110;
        rom_memory[52081] = 3'b110;
        rom_memory[52082] = 3'b110;
        rom_memory[52083] = 3'b110;
        rom_memory[52084] = 3'b110;
        rom_memory[52085] = 3'b110;
        rom_memory[52086] = 3'b110;
        rom_memory[52087] = 3'b110;
        rom_memory[52088] = 3'b111;
        rom_memory[52089] = 3'b111;
        rom_memory[52090] = 3'b111;
        rom_memory[52091] = 3'b111;
        rom_memory[52092] = 3'b110;
        rom_memory[52093] = 3'b110;
        rom_memory[52094] = 3'b110;
        rom_memory[52095] = 3'b110;
        rom_memory[52096] = 3'b110;
        rom_memory[52097] = 3'b110;
        rom_memory[52098] = 3'b100;
        rom_memory[52099] = 3'b100;
        rom_memory[52100] = 3'b100;
        rom_memory[52101] = 3'b100;
        rom_memory[52102] = 3'b100;
        rom_memory[52103] = 3'b100;
        rom_memory[52104] = 3'b100;
        rom_memory[52105] = 3'b100;
        rom_memory[52106] = 3'b100;
        rom_memory[52107] = 3'b100;
        rom_memory[52108] = 3'b100;
        rom_memory[52109] = 3'b100;
        rom_memory[52110] = 3'b110;
        rom_memory[52111] = 3'b110;
        rom_memory[52112] = 3'b110;
        rom_memory[52113] = 3'b110;
        rom_memory[52114] = 3'b110;
        rom_memory[52115] = 3'b111;
        rom_memory[52116] = 3'b111;
        rom_memory[52117] = 3'b111;
        rom_memory[52118] = 3'b111;
        rom_memory[52119] = 3'b111;
        rom_memory[52120] = 3'b111;
        rom_memory[52121] = 3'b111;
        rom_memory[52122] = 3'b111;
        rom_memory[52123] = 3'b110;
        rom_memory[52124] = 3'b110;
        rom_memory[52125] = 3'b110;
        rom_memory[52126] = 3'b110;
        rom_memory[52127] = 3'b111;
        rom_memory[52128] = 3'b111;
        rom_memory[52129] = 3'b110;
        rom_memory[52130] = 3'b000;
        rom_memory[52131] = 3'b000;
        rom_memory[52132] = 3'b100;
        rom_memory[52133] = 3'b110;
        rom_memory[52134] = 3'b111;
        rom_memory[52135] = 3'b111;
        rom_memory[52136] = 3'b111;
        rom_memory[52137] = 3'b111;
        rom_memory[52138] = 3'b111;
        rom_memory[52139] = 3'b111;
        rom_memory[52140] = 3'b111;
        rom_memory[52141] = 3'b110;
        rom_memory[52142] = 3'b110;
        rom_memory[52143] = 3'b110;
        rom_memory[52144] = 3'b110;
        rom_memory[52145] = 3'b000;
        rom_memory[52146] = 3'b000;
        rom_memory[52147] = 3'b000;
        rom_memory[52148] = 3'b111;
        rom_memory[52149] = 3'b111;
        rom_memory[52150] = 3'b110;
        rom_memory[52151] = 3'b110;
        rom_memory[52152] = 3'b110;
        rom_memory[52153] = 3'b100;
        rom_memory[52154] = 3'b100;
        rom_memory[52155] = 3'b100;
        rom_memory[52156] = 3'b110;
        rom_memory[52157] = 3'b110;
        rom_memory[52158] = 3'b100;
        rom_memory[52159] = 3'b110;
        rom_memory[52160] = 3'b110;
        rom_memory[52161] = 3'b110;
        rom_memory[52162] = 3'b110;
        rom_memory[52163] = 3'b111;
        rom_memory[52164] = 3'b111;
        rom_memory[52165] = 3'b111;
        rom_memory[52166] = 3'b111;
        rom_memory[52167] = 3'b111;
        rom_memory[52168] = 3'b111;
        rom_memory[52169] = 3'b111;
        rom_memory[52170] = 3'b111;
        rom_memory[52171] = 3'b111;
        rom_memory[52172] = 3'b111;
        rom_memory[52173] = 3'b111;
        rom_memory[52174] = 3'b110;
        rom_memory[52175] = 3'b111;
        rom_memory[52176] = 3'b111;
        rom_memory[52177] = 3'b110;
        rom_memory[52178] = 3'b110;
        rom_memory[52179] = 3'b110;
        rom_memory[52180] = 3'b110;
        rom_memory[52181] = 3'b110;
        rom_memory[52182] = 3'b110;
        rom_memory[52183] = 3'b110;
        rom_memory[52184] = 3'b110;
        rom_memory[52185] = 3'b100;
        rom_memory[52186] = 3'b100;
        rom_memory[52187] = 3'b100;
        rom_memory[52188] = 3'b100;
        rom_memory[52189] = 3'b101;
        rom_memory[52190] = 3'b111;
        rom_memory[52191] = 3'b100;
        rom_memory[52192] = 3'b100;
        rom_memory[52193] = 3'b100;
        rom_memory[52194] = 3'b000;
        rom_memory[52195] = 3'b000;
        rom_memory[52196] = 3'b000;
        rom_memory[52197] = 3'b000;
        rom_memory[52198] = 3'b000;
        rom_memory[52199] = 3'b100;
        rom_memory[52200] = 3'b111;
        rom_memory[52201] = 3'b111;
        rom_memory[52202] = 3'b111;
        rom_memory[52203] = 3'b111;
        rom_memory[52204] = 3'b111;
        rom_memory[52205] = 3'b111;
        rom_memory[52206] = 3'b110;
        rom_memory[52207] = 3'b110;
        rom_memory[52208] = 3'b110;
        rom_memory[52209] = 3'b110;
        rom_memory[52210] = 3'b110;
        rom_memory[52211] = 3'b110;
        rom_memory[52212] = 3'b110;
        rom_memory[52213] = 3'b110;
        rom_memory[52214] = 3'b110;
        rom_memory[52215] = 3'b110;
        rom_memory[52216] = 3'b110;
        rom_memory[52217] = 3'b110;
        rom_memory[52218] = 3'b110;
        rom_memory[52219] = 3'b110;
        rom_memory[52220] = 3'b110;
        rom_memory[52221] = 3'b110;
        rom_memory[52222] = 3'b110;
        rom_memory[52223] = 3'b110;
        rom_memory[52224] = 3'b110;
        rom_memory[52225] = 3'b110;
        rom_memory[52226] = 3'b110;
        rom_memory[52227] = 3'b110;
        rom_memory[52228] = 3'b110;
        rom_memory[52229] = 3'b110;
        rom_memory[52230] = 3'b110;
        rom_memory[52231] = 3'b110;
        rom_memory[52232] = 3'b110;
        rom_memory[52233] = 3'b110;
        rom_memory[52234] = 3'b110;
        rom_memory[52235] = 3'b110;
        rom_memory[52236] = 3'b110;
        rom_memory[52237] = 3'b110;
        rom_memory[52238] = 3'b110;
        rom_memory[52239] = 3'b111;
        rom_memory[52240] = 3'b111;
        rom_memory[52241] = 3'b111;
        rom_memory[52242] = 3'b111;
        rom_memory[52243] = 3'b111;
        rom_memory[52244] = 3'b111;
        rom_memory[52245] = 3'b111;
        rom_memory[52246] = 3'b111;
        rom_memory[52247] = 3'b111;
        rom_memory[52248] = 3'b111;
        rom_memory[52249] = 3'b111;
        rom_memory[52250] = 3'b111;
        rom_memory[52251] = 3'b111;
        rom_memory[52252] = 3'b111;
        rom_memory[52253] = 3'b111;
        rom_memory[52254] = 3'b111;
        rom_memory[52255] = 3'b111;
        rom_memory[52256] = 3'b111;
        rom_memory[52257] = 3'b111;
        rom_memory[52258] = 3'b111;
        rom_memory[52259] = 3'b111;
        rom_memory[52260] = 3'b111;
        rom_memory[52261] = 3'b111;
        rom_memory[52262] = 3'b111;
        rom_memory[52263] = 3'b111;
        rom_memory[52264] = 3'b111;
        rom_memory[52265] = 3'b111;
        rom_memory[52266] = 3'b111;
        rom_memory[52267] = 3'b111;
        rom_memory[52268] = 3'b111;
        rom_memory[52269] = 3'b111;
        rom_memory[52270] = 3'b111;
        rom_memory[52271] = 3'b111;
        rom_memory[52272] = 3'b111;
        rom_memory[52273] = 3'b111;
        rom_memory[52274] = 3'b111;
        rom_memory[52275] = 3'b111;
        rom_memory[52276] = 3'b111;
        rom_memory[52277] = 3'b111;
        rom_memory[52278] = 3'b111;
        rom_memory[52279] = 3'b111;
        rom_memory[52280] = 3'b111;
        rom_memory[52281] = 3'b111;
        rom_memory[52282] = 3'b111;
        rom_memory[52283] = 3'b111;
        rom_memory[52284] = 3'b111;
        rom_memory[52285] = 3'b111;
        rom_memory[52286] = 3'b111;
        rom_memory[52287] = 3'b111;
        rom_memory[52288] = 3'b111;
        rom_memory[52289] = 3'b111;
        rom_memory[52290] = 3'b111;
        rom_memory[52291] = 3'b111;
        rom_memory[52292] = 3'b111;
        rom_memory[52293] = 3'b111;
        rom_memory[52294] = 3'b111;
        rom_memory[52295] = 3'b111;
        rom_memory[52296] = 3'b111;
        rom_memory[52297] = 3'b111;
        rom_memory[52298] = 3'b111;
        rom_memory[52299] = 3'b111;
        rom_memory[52300] = 3'b111;
        rom_memory[52301] = 3'b111;
        rom_memory[52302] = 3'b111;
        rom_memory[52303] = 3'b111;
        rom_memory[52304] = 3'b111;
        rom_memory[52305] = 3'b111;
        rom_memory[52306] = 3'b111;
        rom_memory[52307] = 3'b111;
        rom_memory[52308] = 3'b111;
        rom_memory[52309] = 3'b111;
        rom_memory[52310] = 3'b111;
        rom_memory[52311] = 3'b111;
        rom_memory[52312] = 3'b111;
        rom_memory[52313] = 3'b111;
        rom_memory[52314] = 3'b111;
        rom_memory[52315] = 3'b111;
        rom_memory[52316] = 3'b111;
        rom_memory[52317] = 3'b111;
        rom_memory[52318] = 3'b111;
        rom_memory[52319] = 3'b111;
        rom_memory[52320] = 3'b110;
        rom_memory[52321] = 3'b110;
        rom_memory[52322] = 3'b110;
        rom_memory[52323] = 3'b110;
        rom_memory[52324] = 3'b110;
        rom_memory[52325] = 3'b110;
        rom_memory[52326] = 3'b110;
        rom_memory[52327] = 3'b110;
        rom_memory[52328] = 3'b110;
        rom_memory[52329] = 3'b110;
        rom_memory[52330] = 3'b110;
        rom_memory[52331] = 3'b110;
        rom_memory[52332] = 3'b110;
        rom_memory[52333] = 3'b110;
        rom_memory[52334] = 3'b110;
        rom_memory[52335] = 3'b110;
        rom_memory[52336] = 3'b110;
        rom_memory[52337] = 3'b110;
        rom_memory[52338] = 3'b110;
        rom_memory[52339] = 3'b100;
        rom_memory[52340] = 3'b100;
        rom_memory[52341] = 3'b100;
        rom_memory[52342] = 3'b100;
        rom_memory[52343] = 3'b100;
        rom_memory[52344] = 3'b100;
        rom_memory[52345] = 3'b100;
        rom_memory[52346] = 3'b100;
        rom_memory[52347] = 3'b100;
        rom_memory[52348] = 3'b100;
        rom_memory[52349] = 3'b100;
        rom_memory[52350] = 3'b110;
        rom_memory[52351] = 3'b110;
        rom_memory[52352] = 3'b110;
        rom_memory[52353] = 3'b110;
        rom_memory[52354] = 3'b110;
        rom_memory[52355] = 3'b111;
        rom_memory[52356] = 3'b111;
        rom_memory[52357] = 3'b111;
        rom_memory[52358] = 3'b111;
        rom_memory[52359] = 3'b111;
        rom_memory[52360] = 3'b111;
        rom_memory[52361] = 3'b111;
        rom_memory[52362] = 3'b111;
        rom_memory[52363] = 3'b111;
        rom_memory[52364] = 3'b111;
        rom_memory[52365] = 3'b111;
        rom_memory[52366] = 3'b110;
        rom_memory[52367] = 3'b111;
        rom_memory[52368] = 3'b111;
        rom_memory[52369] = 3'b111;
        rom_memory[52370] = 3'b100;
        rom_memory[52371] = 3'b000;
        rom_memory[52372] = 3'b111;
        rom_memory[52373] = 3'b111;
        rom_memory[52374] = 3'b111;
        rom_memory[52375] = 3'b111;
        rom_memory[52376] = 3'b111;
        rom_memory[52377] = 3'b111;
        rom_memory[52378] = 3'b111;
        rom_memory[52379] = 3'b111;
        rom_memory[52380] = 3'b111;
        rom_memory[52381] = 3'b110;
        rom_memory[52382] = 3'b110;
        rom_memory[52383] = 3'b110;
        rom_memory[52384] = 3'b110;
        rom_memory[52385] = 3'b000;
        rom_memory[52386] = 3'b000;
        rom_memory[52387] = 3'b000;
        rom_memory[52388] = 3'b110;
        rom_memory[52389] = 3'b110;
        rom_memory[52390] = 3'b100;
        rom_memory[52391] = 3'b110;
        rom_memory[52392] = 3'b110;
        rom_memory[52393] = 3'b100;
        rom_memory[52394] = 3'b100;
        rom_memory[52395] = 3'b110;
        rom_memory[52396] = 3'b111;
        rom_memory[52397] = 3'b111;
        rom_memory[52398] = 3'b111;
        rom_memory[52399] = 3'b111;
        rom_memory[52400] = 3'b110;
        rom_memory[52401] = 3'b111;
        rom_memory[52402] = 3'b111;
        rom_memory[52403] = 3'b111;
        rom_memory[52404] = 3'b111;
        rom_memory[52405] = 3'b111;
        rom_memory[52406] = 3'b111;
        rom_memory[52407] = 3'b111;
        rom_memory[52408] = 3'b111;
        rom_memory[52409] = 3'b111;
        rom_memory[52410] = 3'b111;
        rom_memory[52411] = 3'b110;
        rom_memory[52412] = 3'b110;
        rom_memory[52413] = 3'b110;
        rom_memory[52414] = 3'b110;
        rom_memory[52415] = 3'b110;
        rom_memory[52416] = 3'b110;
        rom_memory[52417] = 3'b110;
        rom_memory[52418] = 3'b110;
        rom_memory[52419] = 3'b110;
        rom_memory[52420] = 3'b110;
        rom_memory[52421] = 3'b110;
        rom_memory[52422] = 3'b110;
        rom_memory[52423] = 3'b000;
        rom_memory[52424] = 3'b000;
        rom_memory[52425] = 3'b000;
        rom_memory[52426] = 3'b000;
        rom_memory[52427] = 3'b100;
        rom_memory[52428] = 3'b100;
        rom_memory[52429] = 3'b100;
        rom_memory[52430] = 3'b100;
        rom_memory[52431] = 3'b100;
        rom_memory[52432] = 3'b100;
        rom_memory[52433] = 3'b100;
        rom_memory[52434] = 3'b000;
        rom_memory[52435] = 3'b000;
        rom_memory[52436] = 3'b000;
        rom_memory[52437] = 3'b000;
        rom_memory[52438] = 3'b000;
        rom_memory[52439] = 3'b000;
        rom_memory[52440] = 3'b100;
        rom_memory[52441] = 3'b111;
        rom_memory[52442] = 3'b111;
        rom_memory[52443] = 3'b111;
        rom_memory[52444] = 3'b111;
        rom_memory[52445] = 3'b111;
        rom_memory[52446] = 3'b111;
        rom_memory[52447] = 3'b110;
        rom_memory[52448] = 3'b110;
        rom_memory[52449] = 3'b110;
        rom_memory[52450] = 3'b110;
        rom_memory[52451] = 3'b110;
        rom_memory[52452] = 3'b110;
        rom_memory[52453] = 3'b110;
        rom_memory[52454] = 3'b110;
        rom_memory[52455] = 3'b110;
        rom_memory[52456] = 3'b110;
        rom_memory[52457] = 3'b110;
        rom_memory[52458] = 3'b110;
        rom_memory[52459] = 3'b110;
        rom_memory[52460] = 3'b110;
        rom_memory[52461] = 3'b110;
        rom_memory[52462] = 3'b110;
        rom_memory[52463] = 3'b110;
        rom_memory[52464] = 3'b110;
        rom_memory[52465] = 3'b110;
        rom_memory[52466] = 3'b110;
        rom_memory[52467] = 3'b110;
        rom_memory[52468] = 3'b110;
        rom_memory[52469] = 3'b110;
        rom_memory[52470] = 3'b110;
        rom_memory[52471] = 3'b110;
        rom_memory[52472] = 3'b110;
        rom_memory[52473] = 3'b110;
        rom_memory[52474] = 3'b110;
        rom_memory[52475] = 3'b110;
        rom_memory[52476] = 3'b110;
        rom_memory[52477] = 3'b110;
        rom_memory[52478] = 3'b110;
        rom_memory[52479] = 3'b111;
        rom_memory[52480] = 3'b111;
        rom_memory[52481] = 3'b111;
        rom_memory[52482] = 3'b111;
        rom_memory[52483] = 3'b111;
        rom_memory[52484] = 3'b111;
        rom_memory[52485] = 3'b111;
        rom_memory[52486] = 3'b111;
        rom_memory[52487] = 3'b111;
        rom_memory[52488] = 3'b111;
        rom_memory[52489] = 3'b111;
        rom_memory[52490] = 3'b111;
        rom_memory[52491] = 3'b111;
        rom_memory[52492] = 3'b111;
        rom_memory[52493] = 3'b111;
        rom_memory[52494] = 3'b111;
        rom_memory[52495] = 3'b111;
        rom_memory[52496] = 3'b111;
        rom_memory[52497] = 3'b111;
        rom_memory[52498] = 3'b111;
        rom_memory[52499] = 3'b111;
        rom_memory[52500] = 3'b111;
        rom_memory[52501] = 3'b111;
        rom_memory[52502] = 3'b111;
        rom_memory[52503] = 3'b111;
        rom_memory[52504] = 3'b111;
        rom_memory[52505] = 3'b111;
        rom_memory[52506] = 3'b111;
        rom_memory[52507] = 3'b111;
        rom_memory[52508] = 3'b111;
        rom_memory[52509] = 3'b111;
        rom_memory[52510] = 3'b111;
        rom_memory[52511] = 3'b111;
        rom_memory[52512] = 3'b111;
        rom_memory[52513] = 3'b111;
        rom_memory[52514] = 3'b111;
        rom_memory[52515] = 3'b111;
        rom_memory[52516] = 3'b111;
        rom_memory[52517] = 3'b111;
        rom_memory[52518] = 3'b111;
        rom_memory[52519] = 3'b111;
        rom_memory[52520] = 3'b111;
        rom_memory[52521] = 3'b111;
        rom_memory[52522] = 3'b111;
        rom_memory[52523] = 3'b111;
        rom_memory[52524] = 3'b111;
        rom_memory[52525] = 3'b111;
        rom_memory[52526] = 3'b111;
        rom_memory[52527] = 3'b111;
        rom_memory[52528] = 3'b111;
        rom_memory[52529] = 3'b111;
        rom_memory[52530] = 3'b111;
        rom_memory[52531] = 3'b111;
        rom_memory[52532] = 3'b111;
        rom_memory[52533] = 3'b111;
        rom_memory[52534] = 3'b111;
        rom_memory[52535] = 3'b111;
        rom_memory[52536] = 3'b111;
        rom_memory[52537] = 3'b111;
        rom_memory[52538] = 3'b111;
        rom_memory[52539] = 3'b111;
        rom_memory[52540] = 3'b111;
        rom_memory[52541] = 3'b111;
        rom_memory[52542] = 3'b111;
        rom_memory[52543] = 3'b111;
        rom_memory[52544] = 3'b111;
        rom_memory[52545] = 3'b111;
        rom_memory[52546] = 3'b111;
        rom_memory[52547] = 3'b111;
        rom_memory[52548] = 3'b111;
        rom_memory[52549] = 3'b111;
        rom_memory[52550] = 3'b111;
        rom_memory[52551] = 3'b111;
        rom_memory[52552] = 3'b111;
        rom_memory[52553] = 3'b111;
        rom_memory[52554] = 3'b111;
        rom_memory[52555] = 3'b111;
        rom_memory[52556] = 3'b111;
        rom_memory[52557] = 3'b111;
        rom_memory[52558] = 3'b111;
        rom_memory[52559] = 3'b111;
        rom_memory[52560] = 3'b110;
        rom_memory[52561] = 3'b110;
        rom_memory[52562] = 3'b110;
        rom_memory[52563] = 3'b110;
        rom_memory[52564] = 3'b110;
        rom_memory[52565] = 3'b110;
        rom_memory[52566] = 3'b110;
        rom_memory[52567] = 3'b110;
        rom_memory[52568] = 3'b110;
        rom_memory[52569] = 3'b110;
        rom_memory[52570] = 3'b110;
        rom_memory[52571] = 3'b110;
        rom_memory[52572] = 3'b110;
        rom_memory[52573] = 3'b110;
        rom_memory[52574] = 3'b110;
        rom_memory[52575] = 3'b110;
        rom_memory[52576] = 3'b110;
        rom_memory[52577] = 3'b110;
        rom_memory[52578] = 3'b110;
        rom_memory[52579] = 3'b100;
        rom_memory[52580] = 3'b100;
        rom_memory[52581] = 3'b100;
        rom_memory[52582] = 3'b100;
        rom_memory[52583] = 3'b100;
        rom_memory[52584] = 3'b100;
        rom_memory[52585] = 3'b100;
        rom_memory[52586] = 3'b100;
        rom_memory[52587] = 3'b100;
        rom_memory[52588] = 3'b100;
        rom_memory[52589] = 3'b100;
        rom_memory[52590] = 3'b110;
        rom_memory[52591] = 3'b110;
        rom_memory[52592] = 3'b110;
        rom_memory[52593] = 3'b110;
        rom_memory[52594] = 3'b110;
        rom_memory[52595] = 3'b111;
        rom_memory[52596] = 3'b111;
        rom_memory[52597] = 3'b111;
        rom_memory[52598] = 3'b111;
        rom_memory[52599] = 3'b111;
        rom_memory[52600] = 3'b111;
        rom_memory[52601] = 3'b111;
        rom_memory[52602] = 3'b111;
        rom_memory[52603] = 3'b111;
        rom_memory[52604] = 3'b111;
        rom_memory[52605] = 3'b111;
        rom_memory[52606] = 3'b110;
        rom_memory[52607] = 3'b111;
        rom_memory[52608] = 3'b111;
        rom_memory[52609] = 3'b111;
        rom_memory[52610] = 3'b111;
        rom_memory[52611] = 3'b100;
        rom_memory[52612] = 3'b100;
        rom_memory[52613] = 3'b111;
        rom_memory[52614] = 3'b111;
        rom_memory[52615] = 3'b111;
        rom_memory[52616] = 3'b111;
        rom_memory[52617] = 3'b111;
        rom_memory[52618] = 3'b111;
        rom_memory[52619] = 3'b111;
        rom_memory[52620] = 3'b111;
        rom_memory[52621] = 3'b110;
        rom_memory[52622] = 3'b110;
        rom_memory[52623] = 3'b110;
        rom_memory[52624] = 3'b110;
        rom_memory[52625] = 3'b000;
        rom_memory[52626] = 3'b000;
        rom_memory[52627] = 3'b000;
        rom_memory[52628] = 3'b000;
        rom_memory[52629] = 3'b110;
        rom_memory[52630] = 3'b100;
        rom_memory[52631] = 3'b100;
        rom_memory[52632] = 3'b100;
        rom_memory[52633] = 3'b110;
        rom_memory[52634] = 3'b111;
        rom_memory[52635] = 3'b111;
        rom_memory[52636] = 3'b111;
        rom_memory[52637] = 3'b111;
        rom_memory[52638] = 3'b111;
        rom_memory[52639] = 3'b111;
        rom_memory[52640] = 3'b111;
        rom_memory[52641] = 3'b111;
        rom_memory[52642] = 3'b111;
        rom_memory[52643] = 3'b111;
        rom_memory[52644] = 3'b111;
        rom_memory[52645] = 3'b111;
        rom_memory[52646] = 3'b111;
        rom_memory[52647] = 3'b111;
        rom_memory[52648] = 3'b111;
        rom_memory[52649] = 3'b110;
        rom_memory[52650] = 3'b110;
        rom_memory[52651] = 3'b110;
        rom_memory[52652] = 3'b110;
        rom_memory[52653] = 3'b110;
        rom_memory[52654] = 3'b110;
        rom_memory[52655] = 3'b110;
        rom_memory[52656] = 3'b110;
        rom_memory[52657] = 3'b110;
        rom_memory[52658] = 3'b110;
        rom_memory[52659] = 3'b110;
        rom_memory[52660] = 3'b100;
        rom_memory[52661] = 3'b000;
        rom_memory[52662] = 3'b000;
        rom_memory[52663] = 3'b000;
        rom_memory[52664] = 3'b000;
        rom_memory[52665] = 3'b000;
        rom_memory[52666] = 3'b000;
        rom_memory[52667] = 3'b100;
        rom_memory[52668] = 3'b100;
        rom_memory[52669] = 3'b100;
        rom_memory[52670] = 3'b100;
        rom_memory[52671] = 3'b100;
        rom_memory[52672] = 3'b100;
        rom_memory[52673] = 3'b100;
        rom_memory[52674] = 3'b100;
        rom_memory[52675] = 3'b000;
        rom_memory[52676] = 3'b000;
        rom_memory[52677] = 3'b000;
        rom_memory[52678] = 3'b000;
        rom_memory[52679] = 3'b000;
        rom_memory[52680] = 3'b100;
        rom_memory[52681] = 3'b101;
        rom_memory[52682] = 3'b111;
        rom_memory[52683] = 3'b111;
        rom_memory[52684] = 3'b111;
        rom_memory[52685] = 3'b111;
        rom_memory[52686] = 3'b111;
        rom_memory[52687] = 3'b110;
        rom_memory[52688] = 3'b110;
        rom_memory[52689] = 3'b110;
        rom_memory[52690] = 3'b110;
        rom_memory[52691] = 3'b110;
        rom_memory[52692] = 3'b110;
        rom_memory[52693] = 3'b110;
        rom_memory[52694] = 3'b110;
        rom_memory[52695] = 3'b110;
        rom_memory[52696] = 3'b110;
        rom_memory[52697] = 3'b110;
        rom_memory[52698] = 3'b110;
        rom_memory[52699] = 3'b110;
        rom_memory[52700] = 3'b110;
        rom_memory[52701] = 3'b110;
        rom_memory[52702] = 3'b110;
        rom_memory[52703] = 3'b110;
        rom_memory[52704] = 3'b110;
        rom_memory[52705] = 3'b110;
        rom_memory[52706] = 3'b110;
        rom_memory[52707] = 3'b110;
        rom_memory[52708] = 3'b110;
        rom_memory[52709] = 3'b110;
        rom_memory[52710] = 3'b110;
        rom_memory[52711] = 3'b110;
        rom_memory[52712] = 3'b110;
        rom_memory[52713] = 3'b110;
        rom_memory[52714] = 3'b110;
        rom_memory[52715] = 3'b110;
        rom_memory[52716] = 3'b110;
        rom_memory[52717] = 3'b110;
        rom_memory[52718] = 3'b111;
        rom_memory[52719] = 3'b111;
        rom_memory[52720] = 3'b111;
        rom_memory[52721] = 3'b111;
        rom_memory[52722] = 3'b111;
        rom_memory[52723] = 3'b111;
        rom_memory[52724] = 3'b111;
        rom_memory[52725] = 3'b111;
        rom_memory[52726] = 3'b111;
        rom_memory[52727] = 3'b111;
        rom_memory[52728] = 3'b111;
        rom_memory[52729] = 3'b111;
        rom_memory[52730] = 3'b111;
        rom_memory[52731] = 3'b111;
        rom_memory[52732] = 3'b111;
        rom_memory[52733] = 3'b111;
        rom_memory[52734] = 3'b111;
        rom_memory[52735] = 3'b111;
        rom_memory[52736] = 3'b111;
        rom_memory[52737] = 3'b111;
        rom_memory[52738] = 3'b111;
        rom_memory[52739] = 3'b111;
        rom_memory[52740] = 3'b111;
        rom_memory[52741] = 3'b111;
        rom_memory[52742] = 3'b111;
        rom_memory[52743] = 3'b111;
        rom_memory[52744] = 3'b111;
        rom_memory[52745] = 3'b111;
        rom_memory[52746] = 3'b111;
        rom_memory[52747] = 3'b111;
        rom_memory[52748] = 3'b111;
        rom_memory[52749] = 3'b111;
        rom_memory[52750] = 3'b111;
        rom_memory[52751] = 3'b111;
        rom_memory[52752] = 3'b111;
        rom_memory[52753] = 3'b111;
        rom_memory[52754] = 3'b111;
        rom_memory[52755] = 3'b111;
        rom_memory[52756] = 3'b111;
        rom_memory[52757] = 3'b111;
        rom_memory[52758] = 3'b111;
        rom_memory[52759] = 3'b111;
        rom_memory[52760] = 3'b111;
        rom_memory[52761] = 3'b111;
        rom_memory[52762] = 3'b111;
        rom_memory[52763] = 3'b111;
        rom_memory[52764] = 3'b111;
        rom_memory[52765] = 3'b111;
        rom_memory[52766] = 3'b111;
        rom_memory[52767] = 3'b111;
        rom_memory[52768] = 3'b111;
        rom_memory[52769] = 3'b111;
        rom_memory[52770] = 3'b111;
        rom_memory[52771] = 3'b111;
        rom_memory[52772] = 3'b111;
        rom_memory[52773] = 3'b111;
        rom_memory[52774] = 3'b111;
        rom_memory[52775] = 3'b111;
        rom_memory[52776] = 3'b111;
        rom_memory[52777] = 3'b111;
        rom_memory[52778] = 3'b111;
        rom_memory[52779] = 3'b111;
        rom_memory[52780] = 3'b111;
        rom_memory[52781] = 3'b111;
        rom_memory[52782] = 3'b111;
        rom_memory[52783] = 3'b111;
        rom_memory[52784] = 3'b111;
        rom_memory[52785] = 3'b111;
        rom_memory[52786] = 3'b111;
        rom_memory[52787] = 3'b111;
        rom_memory[52788] = 3'b111;
        rom_memory[52789] = 3'b111;
        rom_memory[52790] = 3'b111;
        rom_memory[52791] = 3'b111;
        rom_memory[52792] = 3'b111;
        rom_memory[52793] = 3'b111;
        rom_memory[52794] = 3'b111;
        rom_memory[52795] = 3'b111;
        rom_memory[52796] = 3'b111;
        rom_memory[52797] = 3'b111;
        rom_memory[52798] = 3'b111;
        rom_memory[52799] = 3'b111;
    end

    always @(*) begin
        data = rom_memory[addr];
    end
endmodule
